`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.03.2022 17:58:14
// Design Name: 
// Module Name: Note_Displayer
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Note_Displayer(
    input [31:0] freq,
    input CLK100MHZ,
    
    output JC1,JC2,JC3,JC4,JC5,JC6,JC7, JC8
    );
    
    wire [15:0]x;
    wire [15:0]y;
        
    wire frame_begin;
    wire [12:0]pixel_index;
    wire sending_pixels;
    wire sample_pixel;
    wire teststate;
        
    reg [15:0]oled_data; 
    
    my_clock tut4(CLK100MHZ,16,clk6p25m);
    wire clk6p25m;
    wire _20khz_clock;
    my_clock tut3(CLK100MHZ,2499,_20khz_clock);
        
   Oled_Display fnc(clk6p25m, 0, frame_begin, sending_pixels,
        sample_pixel, pixel_index[12:0], oled_data[15:0], JC1, JC2, JC4, JC5, JC6, JC7,
        JC8,teststate);
    
    //letter:(A,0;B,1;C,2;D,3;E,4;F,5;G,6)
    
    
    always @ (posedge CLK100MHZ) begin
    
    if (freq<261 || freq>=2093) //Out_of_Range
    begin
    if (((pixel_index >= 0) && (pixel_index <= 1415)) || ((pixel_index >= 1418) && (pixel_index <= 1465)) || ((pixel_index >= 1471) && (pixel_index <= 1510)) || ((pixel_index >= 1512) && (pixel_index <= 1513)) || ((pixel_index >= 1515) && (pixel_index <= 1560)) || ((pixel_index >= 1563) && (pixel_index <= 1565)) || ((pixel_index >= 1568) && (pixel_index <= 1583)) || ((pixel_index >= 1585) && (pixel_index <= 1605)) || ((pixel_index >= 1608) && (pixel_index <= 1655)) || ((pixel_index >= 1657) && (pixel_index <= 1663)) || ((pixel_index >= 1665) && (pixel_index <= 1679)) || ((pixel_index >= 1681) && (pixel_index <= 1701)) || ((pixel_index >= 1703) && (pixel_index <= 1750)) || ((pixel_index >= 1753) && (pixel_index <= 1759)) || ((pixel_index >= 1762) && (pixel_index <= 1775)) || ((pixel_index >= 1777) && (pixel_index <= 1797)) || ((pixel_index >= 1799) && (pixel_index <= 1846)) || ((pixel_index >= 1848) && (pixel_index <= 1856)) || ((pixel_index >= 1858) && (pixel_index <= 1860)) || ((pixel_index >= 1862) && (pixel_index <= 1866)) || ((pixel_index >= 1868) && (pixel_index <= 1869)) || ((pixel_index >= 1876) && (pixel_index <= 1883)) || ((pixel_index >= 1890) && (pixel_index <= 1892)) || ((pixel_index >= 1898) && (pixel_index <= 1942)) || ((pixel_index >= 1944) && (pixel_index <= 1952)) || ((pixel_index >= 1954) && (pixel_index <= 1956)) || ((pixel_index >= 1958) && (pixel_index <= 1962)) || ((pixel_index >= 1964) && (pixel_index <= 1967)) || ((pixel_index >= 1969) && (pixel_index <= 1978)) || ((pixel_index >= 1981) && (pixel_index <= 1984)) || ((pixel_index >= 1986) && (pixel_index <= 1989)) || ((pixel_index >= 1991) && (pixel_index <= 2038)) || ((pixel_index >= 2040) && (pixel_index <= 2048)) || ((pixel_index >= 2050) && (pixel_index <= 2052)) || ((pixel_index >= 2054) && (pixel_index <= 2058)) || ((pixel_index >= 2060) && (pixel_index <= 2063)) || ((pixel_index >= 2065) && (pixel_index <= 2074)) || ((pixel_index >= 2076) && (pixel_index <= 2080)) || ((pixel_index >= 2083) && (pixel_index <= 2085)) || ((pixel_index >= 2087) && (pixel_index <= 2134)) || ((pixel_index >= 2136) && (pixel_index <= 2144)) || ((pixel_index >= 2146) && (pixel_index <= 2148)) || ((pixel_index >= 2150) && (pixel_index <= 2154)) || ((pixel_index >= 2156) && (pixel_index <= 2159)) || ((pixel_index >= 2161) && (pixel_index <= 2169)) || ((pixel_index >= 2172) && (pixel_index <= 2177)) || ((pixel_index >= 2179) && (pixel_index <= 2181)) || ((pixel_index >= 2183) && (pixel_index <= 2230)) || ((pixel_index >= 2232) && (pixel_index <= 2240)) || ((pixel_index >= 2242) && (pixel_index <= 2244)) || ((pixel_index >= 2246) && (pixel_index <= 2250)) || ((pixel_index >= 2252) && (pixel_index <= 2255)) || ((pixel_index >= 2257) && (pixel_index <= 2265)) || ((pixel_index >= 2268) && (pixel_index <= 2273)) || ((pixel_index >= 2275) && (pixel_index <= 2277)) || ((pixel_index >= 2279) && (pixel_index <= 2326)) || ((pixel_index >= 2328) && (pixel_index <= 2335)) || ((pixel_index >= 2338) && (pixel_index <= 2340)) || ((pixel_index >= 2342) && (pixel_index <= 2346)) || ((pixel_index >= 2348) && (pixel_index <= 2351)) || ((pixel_index >= 2353) && (pixel_index <= 2361)) || ((pixel_index >= 2364) && (pixel_index <= 2369)) || ((pixel_index >= 2371) && (pixel_index <= 2373)) || ((pixel_index >= 2375) && (pixel_index <= 2422)) || ((pixel_index >= 2425) && (pixel_index <= 2431)) || ((pixel_index >= 2433) && (pixel_index <= 2436)) || ((pixel_index >= 2438) && (pixel_index <= 2442)) || ((pixel_index >= 2444) && (pixel_index <= 2447)) || ((pixel_index >= 2449) && (pixel_index <= 2458)) || ((pixel_index >= 2460) && (pixel_index <= 2465)) || ((pixel_index >= 2467) && (pixel_index <= 2469)) || ((pixel_index >= 2471) && (pixel_index <= 2519)) || ((pixel_index >= 2522) && (pixel_index <= 2526)) || ((pixel_index >= 2529) && (pixel_index <= 2532)) || ((pixel_index >= 2534) && (pixel_index <= 2537)) || ((pixel_index >= 2540) && (pixel_index <= 2543)) || ((pixel_index >= 2545) && (pixel_index <= 2554)) || ((pixel_index >= 2556) && (pixel_index <= 2560)) || ((pixel_index >= 2562) && (pixel_index <= 2565)) || ((pixel_index >= 2567) && (pixel_index <= 2616)) || ((pixel_index >= 2624) && (pixel_index <= 2629)) || pixel_index == 2632 || ((pixel_index >= 2636) && (pixel_index <= 2639)) || ((pixel_index >= 2644) && (pixel_index <= 2651)) || ((pixel_index >= 2658) && (pixel_index <= 2661)) || ((pixel_index >= 2663) && (pixel_index <= 2714)) || ((pixel_index >= 2717) && (pixel_index <= 2726)) || ((pixel_index >= 2729) && (pixel_index <= 2737)) || ((pixel_index >= 2739) && (pixel_index <= 2749)) || ((pixel_index >= 2752) && (pixel_index <= 3671)) || ((pixel_index >= 3679) && (pixel_index <= 3767)) || ((pixel_index >= 3770) && (pixel_index <= 3773)) || ((pixel_index >= 3775) && (pixel_index <= 3863)) || ((pixel_index >= 3866) && (pixel_index <= 3869)) || ((pixel_index >= 3872) && (pixel_index <= 3959)) || ((pixel_index >= 3962) && (pixel_index <= 3965)) || ((pixel_index >= 3968) && (pixel_index <= 3971)) || ((pixel_index >= 3976) && (pixel_index <= 3980)) || pixel_index == 3982 || ((pixel_index >= 3987) && (pixel_index <= 3991)) || ((pixel_index >= 3999) && (pixel_index <= 4002)) || ((pixel_index >= 4007) && (pixel_index <= 4055)) || ((pixel_index >= 4058) && (pixel_index <= 4061)) || ((pixel_index >= 4063) && (pixel_index <= 4066)) || ((pixel_index >= 4068) && (pixel_index <= 4071)) || ((pixel_index >= 4073) && (pixel_index <= 4076)) || ((pixel_index >= 4080) && (pixel_index <= 4081)) || ((pixel_index >= 4084) && (pixel_index <= 4086)) || ((pixel_index >= 4089) && (pixel_index <= 4091)) || ((pixel_index >= 4093) && (pixel_index <= 4096)) || ((pixel_index >= 4099) && (pixel_index <= 4101)) || ((pixel_index >= 4104) && (pixel_index <= 4151)) || ((pixel_index >= 4154) && (pixel_index <= 4155)) || ((pixel_index >= 4159) && (pixel_index <= 4167)) || ((pixel_index >= 4169) && (pixel_index <= 4172)) || ((pixel_index >= 4174) && (pixel_index <= 4178)) || ((pixel_index >= 4180) && (pixel_index <= 4182)) || ((pixel_index >= 4184) && (pixel_index <= 4187)) || ((pixel_index >= 4190) && (pixel_index <= 4192)) || ((pixel_index >= 4194) && (pixel_index <= 4198)) || ((pixel_index >= 4200) && (pixel_index <= 4247)) || ((pixel_index >= 4254) && (pixel_index <= 4263)) || ((pixel_index >= 4266) && (pixel_index <= 4268)) || ((pixel_index >= 4270) && (pixel_index <= 4274)) || ((pixel_index >= 4276) && (pixel_index <= 4278)) || ((pixel_index >= 4280) && (pixel_index <= 4284)) || ((pixel_index >= 4286) && (pixel_index <= 4288)) || ((pixel_index >= 4290) && (pixel_index <= 4294)) || ((pixel_index >= 4296) && (pixel_index <= 4343)) || ((pixel_index >= 4346) && (pixel_index <= 4348)) || ((pixel_index >= 4351) && (pixel_index <= 4356)) || ((pixel_index >= 4362) && (pixel_index <= 4364)) || ((pixel_index >= 4366) && (pixel_index <= 4370)) || ((pixel_index >= 4372) && (pixel_index <= 4374)) || ((pixel_index >= 4377) && (pixel_index <= 4379)) || ((pixel_index >= 4382) && (pixel_index <= 4383)) || ((pixel_index >= 4393) && (pixel_index <= 4439)) || ((pixel_index >= 4442) && (pixel_index <= 4445)) || ((pixel_index >= 4447) && (pixel_index <= 4450)) || ((pixel_index >= 4453) && (pixel_index <= 4455)) || ((pixel_index >= 4458) && (pixel_index <= 4460)) || ((pixel_index >= 4462) && (pixel_index <= 4466)) || ((pixel_index >= 4468) && (pixel_index <= 4470)) || ((pixel_index >= 4477) && (pixel_index <= 4479)) || ((pixel_index >= 4482) && (pixel_index <= 4535)) || ((pixel_index >= 4538) && (pixel_index <= 4541)) || ((pixel_index >= 4543) && (pixel_index <= 4546)) || ((pixel_index >= 4548) && (pixel_index <= 4551)) || ((pixel_index >= 4554) && (pixel_index <= 4556)) || ((pixel_index >= 4558) && (pixel_index <= 4562)) || ((pixel_index >= 4564) && (pixel_index <= 4566)) || ((pixel_index >= 4568) && (pixel_index <= 4576)) || ((pixel_index >= 4578) && (pixel_index <= 4631)) || ((pixel_index >= 4634) && (pixel_index <= 4637)) || ((pixel_index >= 4640) && (pixel_index <= 4641)) || ((pixel_index >= 4644) && (pixel_index <= 4647)) || ((pixel_index >= 4650) && (pixel_index <= 4652)) || ((pixel_index >= 4654) && (pixel_index <= 4658)) || ((pixel_index >= 4660) && (pixel_index <= 4662)) || ((pixel_index >= 4664) && (pixel_index <= 4672)) || ((pixel_index >= 4674) && (pixel_index <= 4727)) || ((pixel_index >= 4730) && (pixel_index <= 4734)) || ((pixel_index >= 4736) && (pixel_index <= 4738)) || ((pixel_index >= 4740) && (pixel_index <= 4742)) || ((pixel_index >= 4746) && (pixel_index <= 4748)) || ((pixel_index >= 4750) && (pixel_index <= 4754)) || ((pixel_index >= 4756) && (pixel_index <= 4759)) || ((pixel_index >= 4766) && (pixel_index <= 4768)) || ((pixel_index >= 4771) && (pixel_index <= 4774)) || ((pixel_index >= 4776) && (pixel_index <= 4823)) || ((pixel_index >= 4826) && (pixel_index <= 4830)) || ((pixel_index >= 4833) && (pixel_index <= 4835)) || pixel_index == 4839 || ((pixel_index >= 4842) && (pixel_index <= 4844)) || ((pixel_index >= 4846) && (pixel_index <= 4850)) || ((pixel_index >= 4852) && (pixel_index <= 4854)) || ((pixel_index >= 4856) && (pixel_index <= 4860)) || ((pixel_index >= 4863) && (pixel_index <= 4866)) || ((pixel_index >= 4871) && (pixel_index <= 4950)) || ((pixel_index >= 4952) && (pixel_index <= 4957)) || ((pixel_index >= 4959) && (pixel_index <= 5046)) || ((pixel_index >= 5048) && (pixel_index <= 5052)) || ((pixel_index >= 5055) && (pixel_index <= 5142)) || (pixel_index >= 5150) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1514 || pixel_index == 4087 || pixel_index == 4188 || pixel_index == 4350 || pixel_index == 4832) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2634 || pixel_index == 2642 || pixel_index == 4079 || pixel_index == 4265 || pixel_index == 4361 || pixel_index == 4392 || pixel_index == 4457 || pixel_index == 4553 || pixel_index == 4649 || pixel_index == 4745 || pixel_index == 4841 || pixel_index == 5054) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2751) oled_data = 16'b0101010100001010;
    else oled_data = 0;
    end    
    
    if (freq>=261 && freq<277) //C4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1762)) || ((pixel_index >= 1772) && (pixel_index <= 1788)) || ((pixel_index >= 1793) && (pixel_index <= 1856)) || ((pixel_index >= 1870) && (pixel_index <= 1883)) || ((pixel_index >= 1889) && (pixel_index <= 1951)) || ((pixel_index >= 1956) && (pixel_index <= 1962)) || ((pixel_index >= 1967) && (pixel_index <= 1978)) || ((pixel_index >= 1985) && (pixel_index <= 2046)) || ((pixel_index >= 2051) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2074)) || pixel_index == 2077 || ((pixel_index >= 2081) && (pixel_index <= 2141)) || ((pixel_index >= 2145) && (pixel_index <= 2157)) || ((pixel_index >= 2159) && (pixel_index <= 2169)) || pixel_index == 2173 || ((pixel_index >= 2177) && (pixel_index <= 2237)) || ((pixel_index >= 2241) && (pixel_index <= 2264)) || ((pixel_index >= 2268) && (pixel_index <= 2269)) || ((pixel_index >= 2273) && (pixel_index <= 2332)) || ((pixel_index >= 2336) && (pixel_index <= 2360)) || ((pixel_index >= 2363) && (pixel_index <= 2365)) || ((pixel_index >= 2369) && (pixel_index <= 2428)) || ((pixel_index >= 2432) && (pixel_index <= 2455)) || ((pixel_index >= 2459) && (pixel_index <= 2461)) || ((pixel_index >= 2465) && (pixel_index <= 2524)) || ((pixel_index >= 2527) && (pixel_index <= 2551)) || ((pixel_index >= 2554) && (pixel_index <= 2557)) || ((pixel_index >= 2561) && (pixel_index <= 2619)) || ((pixel_index >= 2623) && (pixel_index <= 2646)) || ((pixel_index >= 2650) && (pixel_index <= 2653)) || ((pixel_index >= 2657) && (pixel_index <= 2715)) || ((pixel_index >= 2719) && (pixel_index <= 2741)) || ((pixel_index >= 2745) && (pixel_index <= 2749)) || ((pixel_index >= 2753) && (pixel_index <= 2811)) || ((pixel_index >= 2815) && (pixel_index <= 2837)) || ((pixel_index >= 2840) && (pixel_index <= 2845)) || ((pixel_index >= 2849) && (pixel_index <= 2907)) || ((pixel_index >= 2911) && (pixel_index <= 2932)) || ((pixel_index >= 2936) && (pixel_index <= 2941)) || ((pixel_index >= 2945) && (pixel_index <= 3003)) || ((pixel_index >= 3007) && (pixel_index <= 3028)) || ((pixel_index >= 3031) && (pixel_index <= 3037)) || ((pixel_index >= 3041) && (pixel_index <= 3099)) || ((pixel_index >= 3103) && (pixel_index <= 3123)) || ((pixel_index >= 3127) && (pixel_index <= 3133)) || ((pixel_index >= 3137) && (pixel_index <= 3195)) || ((pixel_index >= 3199) && (pixel_index <= 3218)) || ((pixel_index >= 3222) && (pixel_index <= 3229)) || ((pixel_index >= 3233) && (pixel_index <= 3291)) || ((pixel_index >= 3295) && (pixel_index <= 3314)) || ((pixel_index >= 3317) && (pixel_index <= 3325)) || ((pixel_index >= 3329) && (pixel_index <= 3387)) || ((pixel_index >= 3391) && (pixel_index <= 3409)) || ((pixel_index >= 3413) && (pixel_index <= 3421)) || ((pixel_index >= 3425) && (pixel_index <= 3483)) || ((pixel_index >= 3487) && (pixel_index <= 3505)) || ((pixel_index >= 3525) && (pixel_index <= 3580)) || ((pixel_index >= 3584) && (pixel_index <= 3601)) || ((pixel_index >= 3621) && (pixel_index <= 3676)) || ((pixel_index >= 3680) && (pixel_index <= 3709)) || ((pixel_index >= 3713) && (pixel_index <= 3773)) || ((pixel_index >= 3777) && (pixel_index <= 3805)) || ((pixel_index >= 3809) && (pixel_index <= 3869)) || ((pixel_index >= 3874) && (pixel_index <= 3885)) || ((pixel_index >= 3887) && (pixel_index <= 3901)) || ((pixel_index >= 3905) && (pixel_index <= 3966)) || ((pixel_index >= 3971) && (pixel_index <= 3979)) || ((pixel_index >= 3983) && (pixel_index <= 3997)) || ((pixel_index >= 4001) && (pixel_index <= 4063)) || ((pixel_index >= 4069) && (pixel_index <= 4073)) || ((pixel_index >= 4079) && (pixel_index <= 4093)) || ((pixel_index >= 4097) && (pixel_index <= 4160)) || ((pixel_index >= 4174) && (pixel_index <= 4189)) || ((pixel_index >= 4193) && (pixel_index <= 4258)) || ((pixel_index >= 4267) && (pixel_index <= 4285)) || (pixel_index >= 4289) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2050 || pixel_index == 2265 || pixel_index == 4173) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=277 && freq<293) //C#4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1389)) || ((pixel_index >= 1392) && (pixel_index <= 1395)) || ((pixel_index >= 1398) && (pixel_index <= 1485)) || ((pixel_index >= 1487) && (pixel_index <= 1491)) || ((pixel_index >= 1493) && (pixel_index <= 1581)) || ((pixel_index >= 1583) && (pixel_index <= 1587)) || ((pixel_index >= 1589) && (pixel_index <= 1676)) || ((pixel_index >= 1679) && (pixel_index <= 1682)) || ((pixel_index >= 1685) && (pixel_index <= 1755)) || ((pixel_index >= 1765) && (pixel_index <= 1772)) || ((pixel_index >= 1775) && (pixel_index <= 1778)) || ((pixel_index >= 1781) && (pixel_index <= 1795)) || ((pixel_index >= 1800) && (pixel_index <= 1849)) || ((pixel_index >= 1863) && (pixel_index <= 1866)) || ((pixel_index >= 1879) && (pixel_index <= 1890)) || ((pixel_index >= 1896) && (pixel_index <= 1944)) || ((pixel_index >= 1949) && (pixel_index <= 1955)) || ((pixel_index >= 1960) && (pixel_index <= 1964)) || ((pixel_index >= 1967) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 1985)) || ((pixel_index >= 1992) && (pixel_index <= 2039)) || ((pixel_index >= 2043) && (pixel_index <= 2053)) || ((pixel_index >= 2056) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2081)) || pixel_index == 2084 || ((pixel_index >= 2088) && (pixel_index <= 2134)) || ((pixel_index >= 2138) && (pixel_index <= 2150)) || ((pixel_index >= 2152) && (pixel_index <= 2156)) || ((pixel_index >= 2159) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2176)) || pixel_index == 2180 || ((pixel_index >= 2184) && (pixel_index <= 2230)) || ((pixel_index >= 2234) && (pixel_index <= 2252)) || ((pixel_index >= 2254) && (pixel_index <= 2258)) || ((pixel_index >= 2260) && (pixel_index <= 2272)) || ((pixel_index >= 2275) && (pixel_index <= 2276)) || ((pixel_index >= 2280) && (pixel_index <= 2325)) || ((pixel_index >= 2329) && (pixel_index <= 2348)) || ((pixel_index >= 2350) && (pixel_index <= 2354)) || ((pixel_index >= 2356) && (pixel_index <= 2367)) || ((pixel_index >= 2371) && (pixel_index <= 2372)) || ((pixel_index >= 2376) && (pixel_index <= 2421)) || ((pixel_index >= 2425) && (pixel_index <= 2441)) || ((pixel_index >= 2454) && (pixel_index <= 2462)) || ((pixel_index >= 2466) && (pixel_index <= 2468)) || ((pixel_index >= 2472) && (pixel_index <= 2516)) || ((pixel_index >= 2520) && (pixel_index <= 2537)) || ((pixel_index >= 2550) && (pixel_index <= 2558)) || ((pixel_index >= 2561) && (pixel_index <= 2564)) || ((pixel_index >= 2568) && (pixel_index <= 2612)) || ((pixel_index >= 2616) && (pixel_index <= 2635)) || ((pixel_index >= 2638) && (pixel_index <= 2641)) || ((pixel_index >= 2644) && (pixel_index <= 2653)) || ((pixel_index >= 2657) && (pixel_index <= 2660)) || ((pixel_index >= 2664) && (pixel_index <= 2708)) || ((pixel_index >= 2712) && (pixel_index <= 2731)) || ((pixel_index >= 2734) && (pixel_index <= 2737)) || ((pixel_index >= 2740) && (pixel_index <= 2749)) || ((pixel_index >= 2752) && (pixel_index <= 2756)) || ((pixel_index >= 2760) && (pixel_index <= 2804)) || ((pixel_index >= 2808) && (pixel_index <= 2827)) || ((pixel_index >= 2830) && (pixel_index <= 2833)) || ((pixel_index >= 2836) && (pixel_index <= 2844)) || ((pixel_index >= 2848) && (pixel_index <= 2852)) || ((pixel_index >= 2856) && (pixel_index <= 2900)) || ((pixel_index >= 2904) && (pixel_index <= 2923)) || ((pixel_index >= 2926) && (pixel_index <= 2929)) || ((pixel_index >= 2932) && (pixel_index <= 2939)) || ((pixel_index >= 2943) && (pixel_index <= 2948)) || ((pixel_index >= 2952) && (pixel_index <= 2996)) || ((pixel_index >= 3000) && (pixel_index <= 3019)) || ((pixel_index >= 3021) && (pixel_index <= 3025)) || ((pixel_index >= 3027) && (pixel_index <= 3035)) || ((pixel_index >= 3038) && (pixel_index <= 3044)) || ((pixel_index >= 3048) && (pixel_index <= 3092)) || ((pixel_index >= 3096) && (pixel_index <= 3130)) || ((pixel_index >= 3134) && (pixel_index <= 3140)) || ((pixel_index >= 3144) && (pixel_index <= 3188)) || ((pixel_index >= 3192) && (pixel_index <= 3226)) || ((pixel_index >= 3229) && (pixel_index <= 3236)) || ((pixel_index >= 3240) && (pixel_index <= 3284)) || ((pixel_index >= 3288) && (pixel_index <= 3321)) || ((pixel_index >= 3325) && (pixel_index <= 3332)) || ((pixel_index >= 3336) && (pixel_index <= 3380)) || ((pixel_index >= 3384) && (pixel_index <= 3416)) || ((pixel_index >= 3420) && (pixel_index <= 3428)) || ((pixel_index >= 3432) && (pixel_index <= 3476)) || ((pixel_index >= 3480) && (pixel_index <= 3512)) || ((pixel_index >= 3532) && (pixel_index <= 3573)) || ((pixel_index >= 3577) && (pixel_index <= 3608)) || ((pixel_index >= 3628) && (pixel_index <= 3669)) || ((pixel_index >= 3673) && (pixel_index <= 3716)) || ((pixel_index >= 3720) && (pixel_index <= 3765)) || ((pixel_index >= 3770) && (pixel_index <= 3812)) || ((pixel_index >= 3816) && (pixel_index <= 3862)) || ((pixel_index >= 3866) && (pixel_index <= 3878)) || ((pixel_index >= 3880) && (pixel_index <= 3908)) || ((pixel_index >= 3912) && (pixel_index <= 3959)) || ((pixel_index >= 3964) && (pixel_index <= 3972)) || ((pixel_index >= 3976) && (pixel_index <= 4004)) || ((pixel_index >= 4008) && (pixel_index <= 4056)) || ((pixel_index >= 4062) && (pixel_index <= 4066)) || ((pixel_index >= 4072) && (pixel_index <= 4100)) || ((pixel_index >= 4104) && (pixel_index <= 4153)) || ((pixel_index >= 4166) && (pixel_index <= 4196)) || ((pixel_index >= 4200) && (pixel_index <= 4251)) || ((pixel_index >= 4260) && (pixel_index <= 4292)) || (pixel_index >= 4296) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1397) oled_data = 16'b0000001010000000;
    else if (pixel_index == 1677 || pixel_index == 2164 || pixel_index == 2370 || pixel_index == 2847) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2931 || pixel_index == 3324) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=293 && freq<311) //D4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1755)) || ((pixel_index >= 1768) && (pixel_index <= 1789)) || ((pixel_index >= 1794) && (pixel_index <= 1851)) || ((pixel_index >= 1866) && (pixel_index <= 1884)) || ((pixel_index >= 1890) && (pixel_index <= 1947)) || ((pixel_index >= 1951) && (pixel_index <= 1957)) || ((pixel_index >= 1964) && (pixel_index <= 1980)) || pixel_index == 1983 || ((pixel_index >= 1986) && (pixel_index <= 2043)) || ((pixel_index >= 2047) && (pixel_index <= 2056)) || ((pixel_index >= 2061) && (pixel_index <= 2075)) || pixel_index == 2079 || ((pixel_index >= 2082) && (pixel_index <= 2139)) || ((pixel_index >= 2143) && (pixel_index <= 2153)) || ((pixel_index >= 2158) && (pixel_index <= 2171)) || ((pixel_index >= 2174) && (pixel_index <= 2175)) || ((pixel_index >= 2178) && (pixel_index <= 2235)) || ((pixel_index >= 2239) && (pixel_index <= 2250)) || ((pixel_index >= 2254) && (pixel_index <= 2266)) || ((pixel_index >= 2270) && (pixel_index <= 2271)) || ((pixel_index >= 2274) && (pixel_index <= 2331)) || ((pixel_index >= 2335) && (pixel_index <= 2347)) || ((pixel_index >= 2351) && (pixel_index <= 2361)) || ((pixel_index >= 2365) && (pixel_index <= 2367)) || ((pixel_index >= 2370) && (pixel_index <= 2427)) || ((pixel_index >= 2431) && (pixel_index <= 2443)) || ((pixel_index >= 2447) && (pixel_index <= 2457)) || ((pixel_index >= 2460) && (pixel_index <= 2463)) || ((pixel_index >= 2466) && (pixel_index <= 2523)) || ((pixel_index >= 2527) && (pixel_index <= 2540)) || ((pixel_index >= 2543) && (pixel_index <= 2552)) || ((pixel_index >= 2556) && (pixel_index <= 2559)) || ((pixel_index >= 2562) && (pixel_index <= 2619)) || ((pixel_index >= 2623) && (pixel_index <= 2636)) || ((pixel_index >= 2640) && (pixel_index <= 2648)) || ((pixel_index >= 2651) && (pixel_index <= 2655)) || ((pixel_index >= 2658) && (pixel_index <= 2715)) || ((pixel_index >= 2719) && (pixel_index <= 2732)) || ((pixel_index >= 2736) && (pixel_index <= 2743)) || ((pixel_index >= 2747) && (pixel_index <= 2751)) || ((pixel_index >= 2754) && (pixel_index <= 2811)) || ((pixel_index >= 2815) && (pixel_index <= 2828)) || ((pixel_index >= 2832) && (pixel_index <= 2838)) || ((pixel_index >= 2842) && (pixel_index <= 2847)) || ((pixel_index >= 2850) && (pixel_index <= 2907)) || ((pixel_index >= 2911) && (pixel_index <= 2924)) || ((pixel_index >= 2928) && (pixel_index <= 2934)) || ((pixel_index >= 2937) && (pixel_index <= 2943)) || ((pixel_index >= 2946) && (pixel_index <= 3003)) || ((pixel_index >= 3007) && (pixel_index <= 3020)) || ((pixel_index >= 3024) && (pixel_index <= 3029)) || ((pixel_index >= 3033) && (pixel_index <= 3039)) || ((pixel_index >= 3042) && (pixel_index <= 3099)) || ((pixel_index >= 3103) && (pixel_index <= 3116)) || ((pixel_index >= 3120) && (pixel_index <= 3125)) || ((pixel_index >= 3128) && (pixel_index <= 3135)) || ((pixel_index >= 3138) && (pixel_index <= 3195)) || ((pixel_index >= 3199) && (pixel_index <= 3212)) || ((pixel_index >= 3216) && (pixel_index <= 3220)) || ((pixel_index >= 3224) && (pixel_index <= 3231)) || ((pixel_index >= 3234) && (pixel_index <= 3291)) || ((pixel_index >= 3295) && (pixel_index <= 3308)) || ((pixel_index >= 3312) && (pixel_index <= 3315)) || ((pixel_index >= 3319) && (pixel_index <= 3327)) || ((pixel_index >= 3330) && (pixel_index <= 3387)) || ((pixel_index >= 3391) && (pixel_index <= 3404)) || ((pixel_index >= 3408) && (pixel_index <= 3411)) || ((pixel_index >= 3414) && (pixel_index <= 3423)) || ((pixel_index >= 3426) && (pixel_index <= 3483)) || ((pixel_index >= 3487) && (pixel_index <= 3499)) || ((pixel_index >= 3503) && (pixel_index <= 3506)) || ((pixel_index >= 3526) && (pixel_index <= 3579)) || ((pixel_index >= 3583) && (pixel_index <= 3595)) || ((pixel_index >= 3599) && (pixel_index <= 3602)) || ((pixel_index >= 3622) && (pixel_index <= 3675)) || ((pixel_index >= 3679) && (pixel_index <= 3691)) || ((pixel_index >= 3695) && (pixel_index <= 3711)) || ((pixel_index >= 3714) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3786)) || ((pixel_index >= 3790) && (pixel_index <= 3807)) || ((pixel_index >= 3810) && (pixel_index <= 3867)) || ((pixel_index >= 3871) && (pixel_index <= 3881)) || ((pixel_index >= 3885) && (pixel_index <= 3903)) || ((pixel_index >= 3906) && (pixel_index <= 3963)) || ((pixel_index >= 3967) && (pixel_index <= 3975)) || ((pixel_index >= 3980) && (pixel_index <= 3999)) || ((pixel_index >= 4002) && (pixel_index <= 4059)) || ((pixel_index >= 4063) && (pixel_index <= 4067)) || ((pixel_index >= 4075) && (pixel_index <= 4095)) || ((pixel_index >= 4098) && (pixel_index <= 4155)) || ((pixel_index >= 4170) && (pixel_index <= 4191)) || ((pixel_index >= 4194) && (pixel_index <= 4251)) || ((pixel_index >= 4263) && (pixel_index <= 4287)) || (pixel_index >= 4290) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 3500 || pixel_index == 4068) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=311 && freq<329) //Eb4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1290)) || ((pixel_index >= 1292) && (pixel_index <= 1386)) || ((pixel_index >= 1388) && (pixel_index <= 1482)) || ((pixel_index >= 1484) && (pixel_index <= 1578)) || ((pixel_index >= 1580) && (pixel_index <= 1674)) || ((pixel_index >= 1676) && (pixel_index <= 1750)) || ((pixel_index >= 1766) && (pixel_index <= 1770)) || ((pixel_index >= 1772) && (pixel_index <= 1794)) || ((pixel_index >= 1799) && (pixel_index <= 1846)) || ((pixel_index >= 1862) && (pixel_index <= 1866)) || ((pixel_index >= 1868) && (pixel_index <= 1869)) || ((pixel_index >= 1875) && (pixel_index <= 1889)) || ((pixel_index >= 1895) && (pixel_index <= 1942)) || ((pixel_index >= 1946) && (pixel_index <= 1962)) || pixel_index == 1964 || ((pixel_index >= 1967) && (pixel_index <= 1969)) || ((pixel_index >= 1972) && (pixel_index <= 1985)) || pixel_index == 1988 || ((pixel_index >= 1991) && (pixel_index <= 2038)) || ((pixel_index >= 2042) && (pixel_index <= 2058)) || ((pixel_index >= 2061) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2080)) || pixel_index == 2084 || ((pixel_index >= 2087) && (pixel_index <= 2134)) || ((pixel_index >= 2138) && (pixel_index <= 2154)) || ((pixel_index >= 2156) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2176)) || ((pixel_index >= 2179) && (pixel_index <= 2180)) || ((pixel_index >= 2183) && (pixel_index <= 2230)) || ((pixel_index >= 2234) && (pixel_index <= 2250)) || ((pixel_index >= 2252) && (pixel_index <= 2259)) || ((pixel_index >= 2261) && (pixel_index <= 2271)) || ((pixel_index >= 2274) && (pixel_index <= 2276)) || ((pixel_index >= 2279) && (pixel_index <= 2326)) || ((pixel_index >= 2330) && (pixel_index <= 2346)) || ((pixel_index >= 2348) && (pixel_index <= 2355)) || ((pixel_index >= 2358) && (pixel_index <= 2366)) || ((pixel_index >= 2370) && (pixel_index <= 2372)) || ((pixel_index >= 2375) && (pixel_index <= 2422)) || ((pixel_index >= 2426) && (pixel_index <= 2442)) || ((pixel_index >= 2444) && (pixel_index <= 2451)) || ((pixel_index >= 2454) && (pixel_index <= 2462)) || ((pixel_index >= 2465) && (pixel_index <= 2468)) || ((pixel_index >= 2471) && (pixel_index <= 2518)) || ((pixel_index >= 2522) && (pixel_index <= 2538)) || ((pixel_index >= 2540) && (pixel_index <= 2547)) || ((pixel_index >= 2549) && (pixel_index <= 2557)) || ((pixel_index >= 2561) && (pixel_index <= 2564)) || ((pixel_index >= 2567) && (pixel_index <= 2614)) || ((pixel_index >= 2618) && (pixel_index <= 2634)) || ((pixel_index >= 2636) && (pixel_index <= 2643)) || ((pixel_index >= 2645) && (pixel_index <= 2652)) || ((pixel_index >= 2656) && (pixel_index <= 2660)) || ((pixel_index >= 2663) && (pixel_index <= 2710)) || ((pixel_index >= 2714) && (pixel_index <= 2730)) || ((pixel_index >= 2732) && (pixel_index <= 2738)) || ((pixel_index >= 2741) && (pixel_index <= 2748)) || ((pixel_index >= 2751) && (pixel_index <= 2756)) || ((pixel_index >= 2759) && (pixel_index <= 2806)) || ((pixel_index >= 2810) && (pixel_index <= 2826)) || ((pixel_index >= 2829) && (pixel_index <= 2834)) || ((pixel_index >= 2837) && (pixel_index <= 2843)) || ((pixel_index >= 2847) && (pixel_index <= 2852)) || ((pixel_index >= 2855) && (pixel_index <= 2902)) || ((pixel_index >= 2916) && (pixel_index <= 2922)) || ((pixel_index >= 2927) && (pixel_index <= 2929)) || ((pixel_index >= 2932) && (pixel_index <= 2939)) || ((pixel_index >= 2942) && (pixel_index <= 2948)) || ((pixel_index >= 2951) && (pixel_index <= 2998)) || ((pixel_index >= 3012) && (pixel_index <= 3018)) || ((pixel_index >= 3020) && (pixel_index <= 3021)) || ((pixel_index >= 3027) && (pixel_index <= 3034)) || ((pixel_index >= 3038) && (pixel_index <= 3044)) || ((pixel_index >= 3047) && (pixel_index <= 3094)) || ((pixel_index >= 3098) && (pixel_index <= 3129)) || ((pixel_index >= 3133) && (pixel_index <= 3140)) || ((pixel_index >= 3143) && (pixel_index <= 3190)) || ((pixel_index >= 3194) && (pixel_index <= 3225)) || ((pixel_index >= 3228) && (pixel_index <= 3236)) || ((pixel_index >= 3239) && (pixel_index <= 3286)) || ((pixel_index >= 3290) && (pixel_index <= 3320)) || ((pixel_index >= 3324) && (pixel_index <= 3332)) || ((pixel_index >= 3335) && (pixel_index <= 3382)) || ((pixel_index >= 3386) && (pixel_index <= 3416)) || ((pixel_index >= 3419) && (pixel_index <= 3428)) || ((pixel_index >= 3431) && (pixel_index <= 3478)) || ((pixel_index >= 3482) && (pixel_index <= 3511)) || ((pixel_index >= 3531) && (pixel_index <= 3574)) || ((pixel_index >= 3578) && (pixel_index <= 3607)) || ((pixel_index >= 3627) && (pixel_index <= 3670)) || ((pixel_index >= 3674) && (pixel_index <= 3716)) || ((pixel_index >= 3719) && (pixel_index <= 3766)) || ((pixel_index >= 3770) && (pixel_index <= 3812)) || ((pixel_index >= 3815) && (pixel_index <= 3862)) || ((pixel_index >= 3866) && (pixel_index <= 3908)) || ((pixel_index >= 3911) && (pixel_index <= 3958)) || ((pixel_index >= 3962) && (pixel_index <= 4004)) || ((pixel_index >= 4007) && (pixel_index <= 4054)) || ((pixel_index >= 4058) && (pixel_index <= 4100)) || ((pixel_index >= 4103) && (pixel_index <= 4150)) || ((pixel_index >= 4166) && (pixel_index <= 4196)) || ((pixel_index >= 4199) && (pixel_index <= 4247)) || ((pixel_index >= 4262) && (pixel_index <= 4292)) || (pixel_index >= 4295) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1765 || pixel_index == 1861 || pixel_index == 2653) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2357 || pixel_index == 3130) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=329 && freq<349) //E4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1758)) || ((pixel_index >= 1773) && (pixel_index <= 1787)) || ((pixel_index >= 1792) && (pixel_index <= 1854)) || ((pixel_index >= 1869) && (pixel_index <= 1882)) || ((pixel_index >= 1888) && (pixel_index <= 1950)) || ((pixel_index >= 1953) && (pixel_index <= 1977)) || ((pixel_index >= 1984) && (pixel_index <= 2046)) || ((pixel_index >= 2049) && (pixel_index <= 2073)) || pixel_index == 2076 || ((pixel_index >= 2080) && (pixel_index <= 2142)) || ((pixel_index >= 2145) && (pixel_index <= 2168)) || pixel_index == 2172 || ((pixel_index >= 2176) && (pixel_index <= 2238)) || ((pixel_index >= 2241) && (pixel_index <= 2264)) || ((pixel_index >= 2267) && (pixel_index <= 2268)) || ((pixel_index >= 2272) && (pixel_index <= 2334)) || ((pixel_index >= 2337) && (pixel_index <= 2359)) || ((pixel_index >= 2362) && (pixel_index <= 2364)) || ((pixel_index >= 2368) && (pixel_index <= 2430)) || ((pixel_index >= 2433) && (pixel_index <= 2454)) || ((pixel_index >= 2458) && (pixel_index <= 2460)) || ((pixel_index >= 2464) && (pixel_index <= 2526)) || ((pixel_index >= 2529) && (pixel_index <= 2550)) || ((pixel_index >= 2553) && (pixel_index <= 2556)) || ((pixel_index >= 2560) && (pixel_index <= 2622)) || ((pixel_index >= 2625) && (pixel_index <= 2645)) || ((pixel_index >= 2649) && (pixel_index <= 2652)) || ((pixel_index >= 2656) && (pixel_index <= 2718)) || ((pixel_index >= 2721) && (pixel_index <= 2740)) || ((pixel_index >= 2744) && (pixel_index <= 2748)) || ((pixel_index >= 2752) && (pixel_index <= 2814)) || ((pixel_index >= 2817) && (pixel_index <= 2836)) || ((pixel_index >= 2839) && (pixel_index <= 2844)) || ((pixel_index >= 2848) && (pixel_index <= 2910)) || ((pixel_index >= 2923) && (pixel_index <= 2931)) || ((pixel_index >= 2935) && (pixel_index <= 2940)) || ((pixel_index >= 2944) && (pixel_index <= 3006)) || ((pixel_index >= 3019) && (pixel_index <= 3027)) || ((pixel_index >= 3030) && (pixel_index <= 3036)) || ((pixel_index >= 3040) && (pixel_index <= 3102)) || ((pixel_index >= 3105) && (pixel_index <= 3122)) || ((pixel_index >= 3126) && (pixel_index <= 3132)) || ((pixel_index >= 3136) && (pixel_index <= 3198)) || ((pixel_index >= 3201) && (pixel_index <= 3217)) || ((pixel_index >= 3221) && (pixel_index <= 3228)) || ((pixel_index >= 3232) && (pixel_index <= 3294)) || ((pixel_index >= 3297) && (pixel_index <= 3313)) || ((pixel_index >= 3316) && (pixel_index <= 3324)) || ((pixel_index >= 3328) && (pixel_index <= 3390)) || ((pixel_index >= 3393) && (pixel_index <= 3408)) || ((pixel_index >= 3412) && (pixel_index <= 3420)) || ((pixel_index >= 3424) && (pixel_index <= 3486)) || ((pixel_index >= 3489) && (pixel_index <= 3504)) || ((pixel_index >= 3524) && (pixel_index <= 3582)) || ((pixel_index >= 3585) && (pixel_index <= 3600)) || ((pixel_index >= 3620) && (pixel_index <= 3678)) || ((pixel_index >= 3681) && (pixel_index <= 3708)) || ((pixel_index >= 3712) && (pixel_index <= 3774)) || ((pixel_index >= 3777) && (pixel_index <= 3804)) || ((pixel_index >= 3808) && (pixel_index <= 3870)) || ((pixel_index >= 3873) && (pixel_index <= 3900)) || ((pixel_index >= 3904) && (pixel_index <= 3966)) || ((pixel_index >= 3969) && (pixel_index <= 3996)) || ((pixel_index >= 4000) && (pixel_index <= 4062)) || ((pixel_index >= 4065) && (pixel_index <= 4092)) || ((pixel_index >= 4096) && (pixel_index <= 4158)) || ((pixel_index >= 4173) && (pixel_index <= 4188)) || ((pixel_index >= 4192) && (pixel_index <= 4254)) || ((pixel_index >= 4269) && (pixel_index <= 4284)) || (pixel_index >= 4288) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2741) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=349 && freq<369) //F4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1758)) || ((pixel_index >= 1773) && (pixel_index <= 1786)) || ((pixel_index >= 1791) && (pixel_index <= 1854)) || ((pixel_index >= 1869) && (pixel_index <= 1881)) || ((pixel_index >= 1887) && (pixel_index <= 1950)) || ((pixel_index >= 1954) && (pixel_index <= 1977)) || pixel_index == 1980 || ((pixel_index >= 1983) && (pixel_index <= 2046)) || ((pixel_index >= 2050) && (pixel_index <= 2072)) || pixel_index == 2076 || ((pixel_index >= 2079) && (pixel_index <= 2142)) || ((pixel_index >= 2146) && (pixel_index <= 2167)) || ((pixel_index >= 2171) && (pixel_index <= 2172)) || ((pixel_index >= 2175) && (pixel_index <= 2238)) || ((pixel_index >= 2242) && (pixel_index <= 2263)) || ((pixel_index >= 2266) && (pixel_index <= 2268)) || ((pixel_index >= 2271) && (pixel_index <= 2334)) || ((pixel_index >= 2338) && (pixel_index <= 2358)) || ((pixel_index >= 2362) && (pixel_index <= 2364)) || ((pixel_index >= 2367) && (pixel_index <= 2430)) || ((pixel_index >= 2434) && (pixel_index <= 2454)) || ((pixel_index >= 2457) && (pixel_index <= 2460)) || ((pixel_index >= 2463) && (pixel_index <= 2526)) || ((pixel_index >= 2530) && (pixel_index <= 2549)) || ((pixel_index >= 2553) && (pixel_index <= 2556)) || ((pixel_index >= 2559) && (pixel_index <= 2622)) || ((pixel_index >= 2626) && (pixel_index <= 2644)) || ((pixel_index >= 2648) && (pixel_index <= 2652)) || ((pixel_index >= 2655) && (pixel_index <= 2718)) || ((pixel_index >= 2722) && (pixel_index <= 2740)) || ((pixel_index >= 2743) && (pixel_index <= 2748)) || ((pixel_index >= 2751) && (pixel_index <= 2814)) || ((pixel_index >= 2818) && (pixel_index <= 2835)) || ((pixel_index >= 2839) && (pixel_index <= 2844)) || ((pixel_index >= 2847) && (pixel_index <= 2910)) || ((pixel_index >= 2924) && (pixel_index <= 2931)) || ((pixel_index >= 2934) && (pixel_index <= 2940)) || ((pixel_index >= 2943) && (pixel_index <= 3006)) || ((pixel_index >= 3020) && (pixel_index <= 3026)) || ((pixel_index >= 3030) && (pixel_index <= 3036)) || ((pixel_index >= 3039) && (pixel_index <= 3102)) || ((pixel_index >= 3116) && (pixel_index <= 3121)) || ((pixel_index >= 3125) && (pixel_index <= 3132)) || ((pixel_index >= 3135) && (pixel_index <= 3198)) || ((pixel_index >= 3202) && (pixel_index <= 3217)) || ((pixel_index >= 3220) && (pixel_index <= 3228)) || ((pixel_index >= 3231) && (pixel_index <= 3294)) || ((pixel_index >= 3298) && (pixel_index <= 3312)) || ((pixel_index >= 3316) && (pixel_index <= 3324)) || ((pixel_index >= 3327) && (pixel_index <= 3390)) || ((pixel_index >= 3394) && (pixel_index <= 3408)) || ((pixel_index >= 3411) && (pixel_index <= 3420)) || ((pixel_index >= 3423) && (pixel_index <= 3486)) || ((pixel_index >= 3490) && (pixel_index <= 3503)) || ((pixel_index >= 3523) && (pixel_index <= 3582)) || ((pixel_index >= 3586) && (pixel_index <= 3599)) || ((pixel_index >= 3619) && (pixel_index <= 3678)) || ((pixel_index >= 3682) && (pixel_index <= 3708)) || ((pixel_index >= 3711) && (pixel_index <= 3774)) || ((pixel_index >= 3778) && (pixel_index <= 3804)) || ((pixel_index >= 3807) && (pixel_index <= 3870)) || ((pixel_index >= 3874) && (pixel_index <= 3900)) || ((pixel_index >= 3903) && (pixel_index <= 3966)) || ((pixel_index >= 3970) && (pixel_index <= 3996)) || ((pixel_index >= 3999) && (pixel_index <= 4062)) || ((pixel_index >= 4066) && (pixel_index <= 4092)) || ((pixel_index >= 4095) && (pixel_index <= 4158)) || ((pixel_index >= 4162) && (pixel_index <= 4188)) || ((pixel_index >= 4191) && (pixel_index <= 4254)) || ((pixel_index >= 4258) && (pixel_index <= 4284)) || (pixel_index >= 4287) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2168) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=369 && freq<391) //F#4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1387)) || ((pixel_index >= 1390) && (pixel_index <= 1393)) || ((pixel_index >= 1396) && (pixel_index <= 1483)) || ((pixel_index >= 1486) && (pixel_index <= 1489)) || ((pixel_index >= 1492) && (pixel_index <= 1579)) || ((pixel_index >= 1582) && (pixel_index <= 1585)) || ((pixel_index >= 1588) && (pixel_index <= 1675)) || ((pixel_index >= 1678) && (pixel_index <= 1681)) || ((pixel_index >= 1684) && (pixel_index <= 1751)) || ((pixel_index >= 1766) && (pixel_index <= 1771)) || ((pixel_index >= 1773) && (pixel_index <= 1777)) || ((pixel_index >= 1779) && (pixel_index <= 1793)) || ((pixel_index >= 1798) && (pixel_index <= 1847)) || ((pixel_index >= 1862) && (pixel_index <= 1864)) || ((pixel_index >= 1878) && (pixel_index <= 1888)) || ((pixel_index >= 1894) && (pixel_index <= 1943)) || ((pixel_index >= 1947) && (pixel_index <= 1962)) || ((pixel_index >= 1965) && (pixel_index <= 1968)) || ((pixel_index >= 1971) && (pixel_index <= 1984)) || pixel_index == 1987 || ((pixel_index >= 1990) && (pixel_index <= 2039)) || ((pixel_index >= 2043) && (pixel_index <= 2058)) || ((pixel_index >= 2061) && (pixel_index <= 2064)) || ((pixel_index >= 2067) && (pixel_index <= 2079)) || pixel_index == 2083 || ((pixel_index >= 2086) && (pixel_index <= 2135)) || ((pixel_index >= 2139) && (pixel_index <= 2154)) || ((pixel_index >= 2157) && (pixel_index <= 2160)) || ((pixel_index >= 2163) && (pixel_index <= 2175)) || ((pixel_index >= 2178) && (pixel_index <= 2179)) || ((pixel_index >= 2182) && (pixel_index <= 2231)) || ((pixel_index >= 2235) && (pixel_index <= 2250)) || ((pixel_index >= 2253) && (pixel_index <= 2256)) || ((pixel_index >= 2259) && (pixel_index <= 2270)) || ((pixel_index >= 2274) && (pixel_index <= 2275)) || ((pixel_index >= 2278) && (pixel_index <= 2327)) || ((pixel_index >= 2331) && (pixel_index <= 2346)) || ((pixel_index >= 2349) && (pixel_index <= 2352)) || ((pixel_index >= 2355) && (pixel_index <= 2365)) || ((pixel_index >= 2369) && (pixel_index <= 2371)) || ((pixel_index >= 2374) && (pixel_index <= 2423)) || ((pixel_index >= 2427) && (pixel_index <= 2440)) || ((pixel_index >= 2453) && (pixel_index <= 2461)) || ((pixel_index >= 2464) && (pixel_index <= 2467)) || ((pixel_index >= 2470) && (pixel_index <= 2519)) || ((pixel_index >= 2523) && (pixel_index <= 2535)) || ((pixel_index >= 2549) && (pixel_index <= 2556)) || ((pixel_index >= 2560) && (pixel_index <= 2563)) || ((pixel_index >= 2566) && (pixel_index <= 2615)) || ((pixel_index >= 2619) && (pixel_index <= 2634)) || ((pixel_index >= 2636) && (pixel_index <= 2640)) || ((pixel_index >= 2642) && (pixel_index <= 2652)) || ((pixel_index >= 2655) && (pixel_index <= 2659)) || ((pixel_index >= 2662) && (pixel_index <= 2711)) || ((pixel_index >= 2715) && (pixel_index <= 2729)) || ((pixel_index >= 2732) && (pixel_index <= 2735)) || ((pixel_index >= 2738) && (pixel_index <= 2747)) || ((pixel_index >= 2751) && (pixel_index <= 2755)) || ((pixel_index >= 2758) && (pixel_index <= 2807)) || ((pixel_index >= 2811) && (pixel_index <= 2825)) || ((pixel_index >= 2828) && (pixel_index <= 2831)) || ((pixel_index >= 2834) && (pixel_index <= 2842)) || ((pixel_index >= 2846) && (pixel_index <= 2851)) || ((pixel_index >= 2854) && (pixel_index <= 2903)) || ((pixel_index >= 2917) && (pixel_index <= 2921)) || ((pixel_index >= 2924) && (pixel_index <= 2927)) || ((pixel_index >= 2930) && (pixel_index <= 2938)) || ((pixel_index >= 2941) && (pixel_index <= 2947)) || ((pixel_index >= 2950) && (pixel_index <= 2999)) || ((pixel_index >= 3013) && (pixel_index <= 3017)) || ((pixel_index >= 3020) && (pixel_index <= 3023)) || ((pixel_index >= 3026) && (pixel_index <= 3033)) || ((pixel_index >= 3037) && (pixel_index <= 3043)) || ((pixel_index >= 3046) && (pixel_index <= 3095)) || ((pixel_index >= 3109) && (pixel_index <= 3129)) || ((pixel_index >= 3132) && (pixel_index <= 3139)) || ((pixel_index >= 3142) && (pixel_index <= 3191)) || ((pixel_index >= 3195) && (pixel_index <= 3224)) || ((pixel_index >= 3228) && (pixel_index <= 3235)) || ((pixel_index >= 3238) && (pixel_index <= 3287)) || ((pixel_index >= 3291) && (pixel_index <= 3319)) || ((pixel_index >= 3323) && (pixel_index <= 3331)) || ((pixel_index >= 3334) && (pixel_index <= 3383)) || ((pixel_index >= 3387) && (pixel_index <= 3415)) || ((pixel_index >= 3418) && (pixel_index <= 3427)) || ((pixel_index >= 3430) && (pixel_index <= 3479)) || ((pixel_index >= 3483) && (pixel_index <= 3510)) || ((pixel_index >= 3530) && (pixel_index <= 3575)) || ((pixel_index >= 3579) && (pixel_index <= 3606)) || ((pixel_index >= 3626) && (pixel_index <= 3671)) || ((pixel_index >= 3675) && (pixel_index <= 3715)) || ((pixel_index >= 3718) && (pixel_index <= 3767)) || ((pixel_index >= 3771) && (pixel_index <= 3811)) || ((pixel_index >= 3814) && (pixel_index <= 3863)) || ((pixel_index >= 3867) && (pixel_index <= 3907)) || ((pixel_index >= 3910) && (pixel_index <= 3959)) || ((pixel_index >= 3963) && (pixel_index <= 4003)) || ((pixel_index >= 4006) && (pixel_index <= 4055)) || ((pixel_index >= 4059) && (pixel_index <= 4099)) || ((pixel_index >= 4102) && (pixel_index <= 4151)) || ((pixel_index >= 4155) && (pixel_index <= 4195)) || ((pixel_index >= 4198) && (pixel_index <= 4247)) || ((pixel_index >= 4251) && (pixel_index <= 4291)) || (pixel_index >= 4294) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1963) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2273 || pixel_index == 2750) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2536 || pixel_index == 3227) oled_data = 16'b1010011110010100;
    else oled_data = 0;
    end
    
    else if (freq>=391 && freq<415) //G4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1761)) || ((pixel_index >= 1772) && (pixel_index <= 1789)) || ((pixel_index >= 1795) && (pixel_index <= 1855)) || ((pixel_index >= 1870) && (pixel_index <= 1885)) || ((pixel_index >= 1891) && (pixel_index <= 1949)) || ((pixel_index >= 1955) && (pixel_index <= 1962)) || ((pixel_index >= 1967) && (pixel_index <= 1980)) || ((pixel_index >= 1987) && (pixel_index <= 2044)) || ((pixel_index >= 2049) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2076)) || pixel_index == 2079 || ((pixel_index >= 2083) && (pixel_index <= 2140)) || ((pixel_index >= 2144) && (pixel_index <= 2171)) || pixel_index == 2175 || ((pixel_index >= 2179) && (pixel_index <= 2235)) || ((pixel_index >= 2239) && (pixel_index <= 2266)) || ((pixel_index >= 2270) && (pixel_index <= 2271)) || ((pixel_index >= 2275) && (pixel_index <= 2330)) || ((pixel_index >= 2334) && (pixel_index <= 2362)) || ((pixel_index >= 2365) && (pixel_index <= 2367)) || ((pixel_index >= 2371) && (pixel_index <= 2426)) || ((pixel_index >= 2430) && (pixel_index <= 2457)) || ((pixel_index >= 2461) && (pixel_index <= 2463)) || ((pixel_index >= 2467) && (pixel_index <= 2522)) || ((pixel_index >= 2525) && (pixel_index <= 2553)) || ((pixel_index >= 2556) && (pixel_index <= 2559)) || ((pixel_index >= 2563) && (pixel_index <= 2617)) || ((pixel_index >= 2621) && (pixel_index <= 2648)) || ((pixel_index >= 2652) && (pixel_index <= 2655)) || ((pixel_index >= 2659) && (pixel_index <= 2713)) || ((pixel_index >= 2717) && (pixel_index <= 2743)) || ((pixel_index >= 2747) && (pixel_index <= 2751)) || ((pixel_index >= 2755) && (pixel_index <= 2809)) || ((pixel_index >= 2813) && (pixel_index <= 2839)) || ((pixel_index >= 2842) && (pixel_index <= 2847)) || ((pixel_index >= 2851) && (pixel_index <= 2905)) || ((pixel_index >= 2909) && (pixel_index <= 2916)) || ((pixel_index >= 2927) && (pixel_index <= 2934)) || ((pixel_index >= 2938) && (pixel_index <= 2943)) || ((pixel_index >= 2947) && (pixel_index <= 3001)) || ((pixel_index >= 3005) && (pixel_index <= 3012)) || ((pixel_index >= 3023) && (pixel_index <= 3030)) || ((pixel_index >= 3033) && (pixel_index <= 3039)) || ((pixel_index >= 3043) && (pixel_index <= 3097)) || ((pixel_index >= 3101) && (pixel_index <= 3108)) || ((pixel_index >= 3119) && (pixel_index <= 3125)) || ((pixel_index >= 3129) && (pixel_index <= 3135)) || ((pixel_index >= 3139) && (pixel_index <= 3193)) || ((pixel_index >= 3197) && (pixel_index <= 3212)) || ((pixel_index >= 3215) && (pixel_index <= 3220)) || ((pixel_index >= 3224) && (pixel_index <= 3231)) || ((pixel_index >= 3235) && (pixel_index <= 3289)) || ((pixel_index >= 3293) && (pixel_index <= 3308)) || ((pixel_index >= 3311) && (pixel_index <= 3316)) || ((pixel_index >= 3319) && (pixel_index <= 3327)) || ((pixel_index >= 3331) && (pixel_index <= 3385)) || ((pixel_index >= 3389) && (pixel_index <= 3404)) || ((pixel_index >= 3407) && (pixel_index <= 3411)) || ((pixel_index >= 3415) && (pixel_index <= 3423)) || ((pixel_index >= 3427) && (pixel_index <= 3482)) || ((pixel_index >= 3486) && (pixel_index <= 3500)) || ((pixel_index >= 3503) && (pixel_index <= 3507)) || ((pixel_index >= 3527) && (pixel_index <= 3578)) || ((pixel_index >= 3582) && (pixel_index <= 3596)) || ((pixel_index >= 3599) && (pixel_index <= 3603)) || ((pixel_index >= 3623) && (pixel_index <= 3674)) || ((pixel_index >= 3679) && (pixel_index <= 3692)) || ((pixel_index >= 3695) && (pixel_index <= 3711)) || ((pixel_index >= 3715) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3788)) || ((pixel_index >= 3791) && (pixel_index <= 3807)) || ((pixel_index >= 3811) && (pixel_index <= 3868)) || ((pixel_index >= 3872) && (pixel_index <= 3884)) || ((pixel_index >= 3887) && (pixel_index <= 3903)) || ((pixel_index >= 3907) && (pixel_index <= 3964)) || ((pixel_index >= 3970) && (pixel_index <= 3979)) || ((pixel_index >= 3983) && (pixel_index <= 3999)) || ((pixel_index >= 4003) && (pixel_index <= 4061)) || ((pixel_index >= 4068) && (pixel_index <= 4073)) || ((pixel_index >= 4079) && (pixel_index <= 4095)) || ((pixel_index >= 4099) && (pixel_index <= 4159)) || ((pixel_index >= 4174) && (pixel_index <= 4191)) || ((pixel_index >= 4195) && (pixel_index <= 4257)) || ((pixel_index >= 4267) && (pixel_index <= 4287)) || (pixel_index >= 4291) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1790) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2267) oled_data = 16'b0000001010000000;
    else if (pixel_index == 2926 || pixel_index == 3485 || pixel_index == 3678) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=415 && freq<440) //Ab4
    begin
    if (((pixel_index >= 0) && (pixel_index <= 1291)) || ((pixel_index >= 1294) && (pixel_index <= 1387)) || ((pixel_index >= 1390) && (pixel_index <= 1483)) || ((pixel_index >= 1486) && (pixel_index <= 1579)) || ((pixel_index >= 1582) && (pixel_index <= 1675)) || ((pixel_index >= 1678) && (pixel_index <= 1755)) || ((pixel_index >= 1759) && (pixel_index <= 1771)) || ((pixel_index >= 1774) && (pixel_index <= 1796)) || ((pixel_index >= 1801) && (pixel_index <= 1851)) || ((pixel_index >= 1856) && (pixel_index <= 1867)) || pixel_index == 1870 || ((pixel_index >= 1877) && (pixel_index <= 1891)) || ((pixel_index >= 1897) && (pixel_index <= 1946)) || ((pixel_index >= 1952) && (pixel_index <= 1963)) || ((pixel_index >= 1968) && (pixel_index <= 1970)) || ((pixel_index >= 1974) && (pixel_index <= 1986)) || ((pixel_index >= 1993) && (pixel_index <= 2042)) || pixel_index == 2045 || ((pixel_index >= 2049) && (pixel_index <= 2059)) || ((pixel_index >= 2063) && (pixel_index <= 2067)) || ((pixel_index >= 2070) && (pixel_index <= 2082)) || pixel_index == 2085 || ((pixel_index >= 2089) && (pixel_index <= 2138)) || pixel_index == 2141 || ((pixel_index >= 2145) && (pixel_index <= 2155)) || ((pixel_index >= 2158) && (pixel_index <= 2164)) || ((pixel_index >= 2167) && (pixel_index <= 2177)) || pixel_index == 2181 || ((pixel_index >= 2185) && (pixel_index <= 2233)) || ((pixel_index >= 2237) && (pixel_index <= 2238)) || ((pixel_index >= 2241) && (pixel_index <= 2251)) || ((pixel_index >= 2254) && (pixel_index <= 2260)) || ((pixel_index >= 2263) && (pixel_index <= 2273)) || ((pixel_index >= 2276) && (pixel_index <= 2277)) || ((pixel_index >= 2281) && (pixel_index <= 2329)) || ((pixel_index >= 2332) && (pixel_index <= 2334)) || ((pixel_index >= 2338) && (pixel_index <= 2347)) || ((pixel_index >= 2350) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2368)) || ((pixel_index >= 2371) && (pixel_index <= 2373)) || ((pixel_index >= 2377) && (pixel_index <= 2424)) || ((pixel_index >= 2428) && (pixel_index <= 2430)) || ((pixel_index >= 2434) && (pixel_index <= 2443)) || ((pixel_index >= 2446) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2463)) || ((pixel_index >= 2467) && (pixel_index <= 2469)) || ((pixel_index >= 2473) && (pixel_index <= 2520)) || ((pixel_index >= 2524) && (pixel_index <= 2527)) || ((pixel_index >= 2530) && (pixel_index <= 2539)) || ((pixel_index >= 2542) && (pixel_index <= 2548)) || ((pixel_index >= 2551) && (pixel_index <= 2559)) || ((pixel_index >= 2562) && (pixel_index <= 2565)) || ((pixel_index >= 2569) && (pixel_index <= 2616)) || ((pixel_index >= 2619) && (pixel_index <= 2623)) || ((pixel_index >= 2627) && (pixel_index <= 2635)) || ((pixel_index >= 2638) && (pixel_index <= 2644)) || ((pixel_index >= 2647) && (pixel_index <= 2654)) || ((pixel_index >= 2658) && (pixel_index <= 2661)) || ((pixel_index >= 2665) && (pixel_index <= 2711)) || ((pixel_index >= 2715) && (pixel_index <= 2719)) || ((pixel_index >= 2723) && (pixel_index <= 2731)) || ((pixel_index >= 2734) && (pixel_index <= 2740)) || ((pixel_index >= 2743) && (pixel_index <= 2749)) || ((pixel_index >= 2753) && (pixel_index <= 2757)) || ((pixel_index >= 2761) && (pixel_index <= 2807)) || ((pixel_index >= 2810) && (pixel_index <= 2816)) || ((pixel_index >= 2820) && (pixel_index <= 2827)) || ((pixel_index >= 2831) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2845)) || ((pixel_index >= 2848) && (pixel_index <= 2853)) || ((pixel_index >= 2857) && (pixel_index <= 2903)) || ((pixel_index >= 2906) && (pixel_index <= 2912)) || ((pixel_index >= 2916) && (pixel_index <= 2923)) || ((pixel_index >= 2928) && (pixel_index <= 2930)) || ((pixel_index >= 2934) && (pixel_index <= 2940)) || ((pixel_index >= 2944) && (pixel_index <= 2949)) || ((pixel_index >= 2953) && (pixel_index <= 2998)) || ((pixel_index >= 3002) && (pixel_index <= 3009)) || ((pixel_index >= 3012) && (pixel_index <= 3019)) || pixel_index == 3022 || ((pixel_index >= 3029) && (pixel_index <= 3036)) || ((pixel_index >= 3039) && (pixel_index <= 3045)) || ((pixel_index >= 3049) && (pixel_index <= 3094)) || ((pixel_index >= 3097) && (pixel_index <= 3105)) || ((pixel_index >= 3109) && (pixel_index <= 3131)) || ((pixel_index >= 3135) && (pixel_index <= 3141)) || ((pixel_index >= 3145) && (pixel_index <= 3190)) || ((pixel_index >= 3193) && (pixel_index <= 3201)) || ((pixel_index >= 3205) && (pixel_index <= 3226)) || ((pixel_index >= 3230) && (pixel_index <= 3237)) || ((pixel_index >= 3241) && (pixel_index <= 3285)) || ((pixel_index >= 3289) && (pixel_index <= 3298)) || ((pixel_index >= 3301) && (pixel_index <= 3322)) || ((pixel_index >= 3325) && (pixel_index <= 3333)) || ((pixel_index >= 3337) && (pixel_index <= 3381)) || ((pixel_index >= 3398) && (pixel_index <= 3417)) || ((pixel_index >= 3421) && (pixel_index <= 3429)) || ((pixel_index >= 3433) && (pixel_index <= 3476)) || ((pixel_index >= 3494) && (pixel_index <= 3513)) || ((pixel_index >= 3533) && (pixel_index <= 3572)) || ((pixel_index >= 3576) && (pixel_index <= 3587)) || ((pixel_index >= 3590) && (pixel_index <= 3609)) || ((pixel_index >= 3629) && (pixel_index <= 3668)) || ((pixel_index >= 3671) && (pixel_index <= 3683)) || ((pixel_index >= 3687) && (pixel_index <= 3717)) || ((pixel_index >= 3721) && (pixel_index <= 3763)) || ((pixel_index >= 3767) && (pixel_index <= 3779)) || ((pixel_index >= 3783) && (pixel_index <= 3813)) || ((pixel_index >= 3817) && (pixel_index <= 3859)) || ((pixel_index >= 3863) && (pixel_index <= 3876)) || ((pixel_index >= 3880) && (pixel_index <= 3909)) || ((pixel_index >= 3913) && (pixel_index <= 3955)) || ((pixel_index >= 3958) && (pixel_index <= 3972)) || ((pixel_index >= 3976) && (pixel_index <= 4005)) || ((pixel_index >= 4009) && (pixel_index <= 4050)) || ((pixel_index >= 4054) && (pixel_index <= 4068)) || ((pixel_index >= 4072) && (pixel_index <= 4101)) || ((pixel_index >= 4105) && (pixel_index <= 4146)) || ((pixel_index >= 4150) && (pixel_index <= 4165)) || ((pixel_index >= 4169) && (pixel_index <= 4197)) || ((pixel_index >= 4201) && (pixel_index <= 4242)) || ((pixel_index >= 4245) && (pixel_index <= 4261)) || ((pixel_index >= 4265) && (pixel_index <= 4293)) || (pixel_index >= 4297) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1971) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2750 || pixel_index == 4069) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2819) oled_data = 16'b0101010100001010;
    else oled_data = 0;
    end
    
    else if (freq>=440 && freq<466) //A4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1762)) || ((pixel_index >= 1767) && (pixel_index <= 1788)) || ((pixel_index >= 1793) && (pixel_index <= 1858)) || ((pixel_index >= 1863) && (pixel_index <= 1884)) || ((pixel_index >= 1889) && (pixel_index <= 1954)) || ((pixel_index >= 1960) && (pixel_index <= 1979)) || pixel_index == 1982 || ((pixel_index >= 1985) && (pixel_index <= 2049)) || ((pixel_index >= 2056) && (pixel_index <= 2074)) || pixel_index == 2078 || ((pixel_index >= 2081) && (pixel_index <= 2145)) || ((pixel_index >= 2148) && (pixel_index <= 2149)) || ((pixel_index >= 2152) && (pixel_index <= 2170)) || ((pixel_index >= 2173) && (pixel_index <= 2174)) || ((pixel_index >= 2177) && (pixel_index <= 2241)) || ((pixel_index >= 2244) && (pixel_index <= 2245)) || ((pixel_index >= 2249) && (pixel_index <= 2265)) || ((pixel_index >= 2269) && (pixel_index <= 2270)) || ((pixel_index >= 2273) && (pixel_index <= 2336)) || ((pixel_index >= 2340) && (pixel_index <= 2341)) || ((pixel_index >= 2345) && (pixel_index <= 2360)) || ((pixel_index >= 2364) && (pixel_index <= 2366)) || ((pixel_index >= 2369) && (pixel_index <= 2432)) || ((pixel_index >= 2435) && (pixel_index <= 2438)) || ((pixel_index >= 2441) && (pixel_index <= 2456)) || ((pixel_index >= 2459) && (pixel_index <= 2462)) || ((pixel_index >= 2465) && (pixel_index <= 2527)) || ((pixel_index >= 2531) && (pixel_index <= 2534)) || ((pixel_index >= 2538) && (pixel_index <= 2551)) || ((pixel_index >= 2555) && (pixel_index <= 2558)) || ((pixel_index >= 2561) && (pixel_index <= 2623)) || ((pixel_index >= 2627) && (pixel_index <= 2630)) || ((pixel_index >= 2634) && (pixel_index <= 2647)) || ((pixel_index >= 2650) && (pixel_index <= 2654)) || ((pixel_index >= 2657) && (pixel_index <= 2719)) || ((pixel_index >= 2722) && (pixel_index <= 2727)) || ((pixel_index >= 2731) && (pixel_index <= 2742)) || ((pixel_index >= 2746) && (pixel_index <= 2750)) || ((pixel_index >= 2753) && (pixel_index <= 2814)) || ((pixel_index >= 2818) && (pixel_index <= 2823)) || ((pixel_index >= 2827) && (pixel_index <= 2837)) || ((pixel_index >= 2841) && (pixel_index <= 2846)) || ((pixel_index >= 2849) && (pixel_index <= 2910)) || ((pixel_index >= 2914) && (pixel_index <= 2920)) || ((pixel_index >= 2923) && (pixel_index <= 2933)) || ((pixel_index >= 2936) && (pixel_index <= 2942)) || ((pixel_index >= 2945) && (pixel_index <= 3006)) || ((pixel_index >= 3009) && (pixel_index <= 3016)) || ((pixel_index >= 3020) && (pixel_index <= 3028)) || ((pixel_index >= 3032) && (pixel_index <= 3038)) || ((pixel_index >= 3041) && (pixel_index <= 3101)) || ((pixel_index >= 3105) && (pixel_index <= 3112)) || ((pixel_index >= 3116) && (pixel_index <= 3124)) || ((pixel_index >= 3127) && (pixel_index <= 3134)) || ((pixel_index >= 3137) && (pixel_index <= 3197)) || ((pixel_index >= 3201) && (pixel_index <= 3209)) || ((pixel_index >= 3212) && (pixel_index <= 3219)) || ((pixel_index >= 3223) && (pixel_index <= 3230)) || ((pixel_index >= 3233) && (pixel_index <= 3293)) || ((pixel_index >= 3296) && (pixel_index <= 3305)) || ((pixel_index >= 3309) && (pixel_index <= 3314)) || ((pixel_index >= 3318) && (pixel_index <= 3326)) || ((pixel_index >= 3329) && (pixel_index <= 3388)) || ((pixel_index >= 3405) && (pixel_index <= 3410)) || ((pixel_index >= 3413) && (pixel_index <= 3422)) || ((pixel_index >= 3425) && (pixel_index <= 3484)) || ((pixel_index >= 3501) && (pixel_index <= 3505)) || ((pixel_index >= 3525) && (pixel_index <= 3579)) || ((pixel_index >= 3583) && (pixel_index <= 3594)) || ((pixel_index >= 3598) && (pixel_index <= 3601)) || ((pixel_index >= 3621) && (pixel_index <= 3675)) || ((pixel_index >= 3679) && (pixel_index <= 3690)) || ((pixel_index >= 3694) && (pixel_index <= 3710)) || ((pixel_index >= 3713) && (pixel_index <= 3771)) || ((pixel_index >= 3774) && (pixel_index <= 3787)) || ((pixel_index >= 3791) && (pixel_index <= 3806)) || ((pixel_index >= 3809) && (pixel_index <= 3866)) || ((pixel_index >= 3870) && (pixel_index <= 3883)) || ((pixel_index >= 3887) && (pixel_index <= 3902)) || ((pixel_index >= 3905) && (pixel_index <= 3962)) || ((pixel_index >= 3966) && (pixel_index <= 3980)) || ((pixel_index >= 3983) && (pixel_index <= 3998)) || ((pixel_index >= 4001) && (pixel_index <= 4058)) || ((pixel_index >= 4061) && (pixel_index <= 4076)) || ((pixel_index >= 4080) && (pixel_index <= 4094)) || ((pixel_index >= 4097) && (pixel_index <= 4153)) || ((pixel_index >= 4157) && (pixel_index <= 4172)) || ((pixel_index >= 4176) && (pixel_index <= 4190)) || ((pixel_index >= 4193) && (pixel_index <= 4249)) || ((pixel_index >= 4253) && (pixel_index <= 4269)) || ((pixel_index >= 4272) && (pixel_index <= 4286)) || (pixel_index >= 4289) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2361 || pixel_index == 2528 || pixel_index == 2631 || pixel_index == 3200) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=466 && freq<493) //Bb4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1290)) || ((pixel_index >= 1293) && (pixel_index <= 1386)) || ((pixel_index >= 1389) && (pixel_index <= 1482)) || ((pixel_index >= 1485) && (pixel_index <= 1578)) || ((pixel_index >= 1581) && (pixel_index <= 1674)) || ((pixel_index >= 1677) && (pixel_index <= 1749)) || ((pixel_index >= 1762) && (pixel_index <= 1770)) || ((pixel_index >= 1773) && (pixel_index <= 1795)) || ((pixel_index >= 1800) && (pixel_index <= 1845)) || ((pixel_index >= 1859) && (pixel_index <= 1866)) || ((pixel_index >= 1869) && (pixel_index <= 1870)) || ((pixel_index >= 1876) && (pixel_index <= 1890)) || ((pixel_index >= 1896) && (pixel_index <= 1941)) || ((pixel_index >= 1945) && (pixel_index <= 1951)) || ((pixel_index >= 1956) && (pixel_index <= 1962)) || ((pixel_index >= 1968) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 1986)) || pixel_index == 1989 || ((pixel_index >= 1992) && (pixel_index <= 2037)) || ((pixel_index >= 2041) && (pixel_index <= 2048)) || ((pixel_index >= 2053) && (pixel_index <= 2058)) || ((pixel_index >= 2062) && (pixel_index <= 2067)) || ((pixel_index >= 2070) && (pixel_index <= 2081)) || pixel_index == 2085 || ((pixel_index >= 2088) && (pixel_index <= 2133)) || ((pixel_index >= 2137) && (pixel_index <= 2145)) || ((pixel_index >= 2149) && (pixel_index <= 2154)) || ((pixel_index >= 2157) && (pixel_index <= 2163)) || ((pixel_index >= 2166) && (pixel_index <= 2177)) || ((pixel_index >= 2180) && (pixel_index <= 2181)) || ((pixel_index >= 2184) && (pixel_index <= 2229)) || ((pixel_index >= 2233) && (pixel_index <= 2241)) || ((pixel_index >= 2245) && (pixel_index <= 2250)) || ((pixel_index >= 2253) && (pixel_index <= 2260)) || ((pixel_index >= 2262) && (pixel_index <= 2272)) || ((pixel_index >= 2275) && (pixel_index <= 2277)) || ((pixel_index >= 2280) && (pixel_index <= 2325)) || ((pixel_index >= 2329) && (pixel_index <= 2338)) || ((pixel_index >= 2341) && (pixel_index <= 2346)) || ((pixel_index >= 2349) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2367)) || ((pixel_index >= 2371) && (pixel_index <= 2373)) || ((pixel_index >= 2376) && (pixel_index <= 2421)) || ((pixel_index >= 2425) && (pixel_index <= 2434)) || ((pixel_index >= 2437) && (pixel_index <= 2442)) || ((pixel_index >= 2445) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2463)) || ((pixel_index >= 2466) && (pixel_index <= 2469)) || ((pixel_index >= 2472) && (pixel_index <= 2517)) || ((pixel_index >= 2521) && (pixel_index <= 2529)) || ((pixel_index >= 2533) && (pixel_index <= 2538)) || ((pixel_index >= 2541) && (pixel_index <= 2548)) || ((pixel_index >= 2550) && (pixel_index <= 2558)) || ((pixel_index >= 2562) && (pixel_index <= 2565)) || ((pixel_index >= 2568) && (pixel_index <= 2613)) || ((pixel_index >= 2617) && (pixel_index <= 2625)) || ((pixel_index >= 2629) && (pixel_index <= 2634)) || ((pixel_index >= 2637) && (pixel_index <= 2644)) || ((pixel_index >= 2646) && (pixel_index <= 2653)) || ((pixel_index >= 2657) && (pixel_index <= 2661)) || ((pixel_index >= 2664) && (pixel_index <= 2709)) || ((pixel_index >= 2713) && (pixel_index <= 2720)) || ((pixel_index >= 2724) && (pixel_index <= 2730)) || ((pixel_index >= 2733) && (pixel_index <= 2739)) || ((pixel_index >= 2742) && (pixel_index <= 2749)) || ((pixel_index >= 2752) && (pixel_index <= 2757)) || ((pixel_index >= 2760) && (pixel_index <= 2805)) || ((pixel_index >= 2809) && (pixel_index <= 2815)) || ((pixel_index >= 2819) && (pixel_index <= 2826)) || ((pixel_index >= 2830) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2844)) || ((pixel_index >= 2848) && (pixel_index <= 2853)) || ((pixel_index >= 2856) && (pixel_index <= 2901)) || ((pixel_index >= 2914) && (pixel_index <= 2922)) || ((pixel_index >= 2928) && (pixel_index <= 2930)) || ((pixel_index >= 2933) && (pixel_index <= 2940)) || ((pixel_index >= 2943) && (pixel_index <= 2949)) || ((pixel_index >= 2952) && (pixel_index <= 2997)) || ((pixel_index >= 3012) && (pixel_index <= 3018)) || ((pixel_index >= 3021) && (pixel_index <= 3022)) || ((pixel_index >= 3028) && (pixel_index <= 3035)) || ((pixel_index >= 3039) && (pixel_index <= 3045)) || ((pixel_index >= 3048) && (pixel_index <= 3093)) || ((pixel_index >= 3097) && (pixel_index <= 3104)) || ((pixel_index >= 3109) && (pixel_index <= 3130)) || ((pixel_index >= 3134) && (pixel_index <= 3141)) || ((pixel_index >= 3144) && (pixel_index <= 3189)) || ((pixel_index >= 3193) && (pixel_index <= 3202)) || ((pixel_index >= 3206) && (pixel_index <= 3226)) || ((pixel_index >= 3229) && (pixel_index <= 3237)) || ((pixel_index >= 3240) && (pixel_index <= 3285)) || ((pixel_index >= 3289) && (pixel_index <= 3299)) || ((pixel_index >= 3303) && (pixel_index <= 3321)) || ((pixel_index >= 3325) && (pixel_index <= 3333)) || ((pixel_index >= 3336) && (pixel_index <= 3381)) || ((pixel_index >= 3385) && (pixel_index <= 3395)) || ((pixel_index >= 3399) && (pixel_index <= 3417)) || ((pixel_index >= 3420) && (pixel_index <= 3429)) || ((pixel_index >= 3432) && (pixel_index <= 3477)) || ((pixel_index >= 3481) && (pixel_index <= 3491)) || ((pixel_index >= 3495) && (pixel_index <= 3512)) || ((pixel_index >= 3532) && (pixel_index <= 3573)) || ((pixel_index >= 3577) && (pixel_index <= 3587)) || ((pixel_index >= 3591) && (pixel_index <= 3608)) || ((pixel_index >= 3628) && (pixel_index <= 3669)) || ((pixel_index >= 3673) && (pixel_index <= 3683)) || ((pixel_index >= 3687) && (pixel_index <= 3717)) || ((pixel_index >= 3720) && (pixel_index <= 3765)) || ((pixel_index >= 3769) && (pixel_index <= 3779)) || ((pixel_index >= 3783) && (pixel_index <= 3813)) || ((pixel_index >= 3816) && (pixel_index <= 3861)) || ((pixel_index >= 3865) && (pixel_index <= 3874)) || ((pixel_index >= 3878) && (pixel_index <= 3909)) || ((pixel_index >= 3912) && (pixel_index <= 3957)) || ((pixel_index >= 3961) && (pixel_index <= 3969)) || ((pixel_index >= 3974) && (pixel_index <= 4005)) || ((pixel_index >= 4008) && (pixel_index <= 4053)) || ((pixel_index >= 4057) && (pixel_index <= 4063)) || ((pixel_index >= 4069) && (pixel_index <= 4101)) || ((pixel_index >= 4104) && (pixel_index <= 4149)) || ((pixel_index >= 4164) && (pixel_index <= 4197)) || ((pixel_index >= 4200) && (pixel_index <= 4246)) || ((pixel_index >= 4258) && (pixel_index <= 4293)) || (pixel_index >= 4296) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1291 || pixel_index == 1387 || pixel_index == 1483 || pixel_index == 1579 || pixel_index == 1675 || pixel_index == 1771 || pixel_index == 1867 || pixel_index == 1963 || pixel_index == 1965 || pixel_index == 2059 || pixel_index == 2155 || pixel_index == 2251 || pixel_index == 2347 || pixel_index == 2358 || pixel_index == 2443 || pixel_index == 2539 || pixel_index == 2635 || pixel_index == 2731 || pixel_index == 2827 || pixel_index == 2923 || pixel_index == 3019) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2049 || pixel_index == 2242 || pixel_index == 2654) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=493 && freq<523) //B4
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1757)) || ((pixel_index >= 1769) && (pixel_index <= 1788)) || ((pixel_index >= 1793) && (pixel_index <= 1853)) || ((pixel_index >= 1867) && (pixel_index <= 1883)) || ((pixel_index >= 1889) && (pixel_index <= 1949)) || ((pixel_index >= 1952) && (pixel_index <= 1958)) || ((pixel_index >= 1964) && (pixel_index <= 1978)) || ((pixel_index >= 1985) && (pixel_index <= 2045)) || ((pixel_index >= 2048) && (pixel_index <= 2056)) || ((pixel_index >= 2060) && (pixel_index <= 2074)) || pixel_index == 2077 || ((pixel_index >= 2081) && (pixel_index <= 2141)) || ((pixel_index >= 2144) && (pixel_index <= 2153)) || ((pixel_index >= 2157) && (pixel_index <= 2169)) || pixel_index == 2173 || ((pixel_index >= 2177) && (pixel_index <= 2237)) || ((pixel_index >= 2240) && (pixel_index <= 2249)) || ((pixel_index >= 2253) && (pixel_index <= 2264)) || ((pixel_index >= 2268) && (pixel_index <= 2269)) || ((pixel_index >= 2273) && (pixel_index <= 2333)) || ((pixel_index >= 2336) && (pixel_index <= 2345)) || ((pixel_index >= 2349) && (pixel_index <= 2360)) || ((pixel_index >= 2363) && (pixel_index <= 2365)) || ((pixel_index >= 2369) && (pixel_index <= 2429)) || ((pixel_index >= 2432) && (pixel_index <= 2441)) || ((pixel_index >= 2445) && (pixel_index <= 2455)) || ((pixel_index >= 2459) && (pixel_index <= 2461)) || ((pixel_index >= 2465) && (pixel_index <= 2525)) || ((pixel_index >= 2528) && (pixel_index <= 2537)) || ((pixel_index >= 2541) && (pixel_index <= 2551)) || ((pixel_index >= 2554) && (pixel_index <= 2557)) || ((pixel_index >= 2561) && (pixel_index <= 2621)) || ((pixel_index >= 2624) && (pixel_index <= 2632)) || ((pixel_index >= 2636) && (pixel_index <= 2646)) || ((pixel_index >= 2650) && (pixel_index <= 2653)) || ((pixel_index >= 2657) && (pixel_index <= 2717)) || ((pixel_index >= 2720) && (pixel_index <= 2728)) || ((pixel_index >= 2732) && (pixel_index <= 2741)) || ((pixel_index >= 2745) && (pixel_index <= 2749)) || ((pixel_index >= 2753) && (pixel_index <= 2813)) || ((pixel_index >= 2816) && (pixel_index <= 2822)) || ((pixel_index >= 2827) && (pixel_index <= 2837)) || ((pixel_index >= 2840) && (pixel_index <= 2845)) || ((pixel_index >= 2849) && (pixel_index <= 2909)) || ((pixel_index >= 2921) && (pixel_index <= 2932)) || ((pixel_index >= 2936) && (pixel_index <= 2941)) || ((pixel_index >= 2945) && (pixel_index <= 3005)) || ((pixel_index >= 3020) && (pixel_index <= 3028)) || ((pixel_index >= 3031) && (pixel_index <= 3037)) || ((pixel_index >= 3041) && (pixel_index <= 3101)) || ((pixel_index >= 3104) && (pixel_index <= 3111)) || ((pixel_index >= 3117) && (pixel_index <= 3123)) || ((pixel_index >= 3127) && (pixel_index <= 3133)) || ((pixel_index >= 3137) && (pixel_index <= 3197)) || ((pixel_index >= 3200) && (pixel_index <= 3209)) || ((pixel_index >= 3214) && (pixel_index <= 3218)) || ((pixel_index >= 3222) && (pixel_index <= 3229)) || ((pixel_index >= 3233) && (pixel_index <= 3293)) || ((pixel_index >= 3296) && (pixel_index <= 3306)) || ((pixel_index >= 3310) && (pixel_index <= 3314)) || ((pixel_index >= 3317) && (pixel_index <= 3325)) || ((pixel_index >= 3329) && (pixel_index <= 3389)) || ((pixel_index >= 3392) && (pixel_index <= 3402)) || ((pixel_index >= 3406) && (pixel_index <= 3409)) || ((pixel_index >= 3413) && (pixel_index <= 3421)) || ((pixel_index >= 3425) && (pixel_index <= 3485)) || ((pixel_index >= 3488) && (pixel_index <= 3499)) || ((pixel_index >= 3503) && (pixel_index <= 3505)) || ((pixel_index >= 3525) && (pixel_index <= 3581)) || ((pixel_index >= 3584) && (pixel_index <= 3595)) || ((pixel_index >= 3599) && (pixel_index <= 3601)) || ((pixel_index >= 3621) && (pixel_index <= 3677)) || ((pixel_index >= 3680) && (pixel_index <= 3691)) || ((pixel_index >= 3694) && (pixel_index <= 3709)) || ((pixel_index >= 3713) && (pixel_index <= 3773)) || ((pixel_index >= 3776) && (pixel_index <= 3786)) || ((pixel_index >= 3790) && (pixel_index <= 3805)) || ((pixel_index >= 3809) && (pixel_index <= 3869)) || ((pixel_index >= 3872) && (pixel_index <= 3882)) || ((pixel_index >= 3886) && (pixel_index <= 3901)) || ((pixel_index >= 3905) && (pixel_index <= 3965)) || ((pixel_index >= 3968) && (pixel_index <= 3977)) || ((pixel_index >= 3981) && (pixel_index <= 3997)) || ((pixel_index >= 4001) && (pixel_index <= 4061)) || ((pixel_index >= 4064) && (pixel_index <= 4070)) || ((pixel_index >= 4077) && (pixel_index <= 4093)) || ((pixel_index >= 4097) && (pixel_index <= 4157)) || ((pixel_index >= 4171) && (pixel_index <= 4189)) || ((pixel_index >= 4193) && (pixel_index <= 4253)) || ((pixel_index >= 4265) && (pixel_index <= 4285)) || (pixel_index >= 4289) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2156 || pixel_index == 3403 || pixel_index == 3598) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2265 || pixel_index == 3213 || pixel_index == 3502) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=523 && freq<554) //C5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1762)) || ((pixel_index >= 1772) && (pixel_index <= 1779)) || ((pixel_index >= 1794) && (pixel_index <= 1856)) || ((pixel_index >= 1870) && (pixel_index <= 1875)) || ((pixel_index >= 1890) && (pixel_index <= 1951)) || ((pixel_index >= 1956) && (pixel_index <= 1962)) || ((pixel_index >= 1967) && (pixel_index <= 1971)) || ((pixel_index >= 1975) && (pixel_index <= 2046)) || ((pixel_index >= 2051) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2067)) || ((pixel_index >= 2071) && (pixel_index <= 2141)) || ((pixel_index >= 2145) && (pixel_index <= 2157)) || ((pixel_index >= 2159) && (pixel_index <= 2163)) || ((pixel_index >= 2167) && (pixel_index <= 2237)) || ((pixel_index >= 2241) && (pixel_index <= 2259)) || ((pixel_index >= 2263) && (pixel_index <= 2332)) || ((pixel_index >= 2336) && (pixel_index <= 2355)) || ((pixel_index >= 2359) && (pixel_index <= 2428)) || ((pixel_index >= 2432) && (pixel_index <= 2451)) || ((pixel_index >= 2455) && (pixel_index <= 2524)) || ((pixel_index >= 2527) && (pixel_index <= 2547)) || ((pixel_index >= 2551) && (pixel_index <= 2619)) || ((pixel_index >= 2623) && (pixel_index <= 2643)) || ((pixel_index >= 2647) && (pixel_index <= 2715)) || ((pixel_index >= 2719) && (pixel_index <= 2739)) || ((pixel_index >= 2743) && (pixel_index <= 2811)) || ((pixel_index >= 2815) && (pixel_index <= 2835)) || ((pixel_index >= 2847) && (pixel_index <= 2907)) || ((pixel_index >= 2911) && (pixel_index <= 2931)) || ((pixel_index >= 2945) && (pixel_index <= 3003)) || ((pixel_index >= 3007) && (pixel_index <= 3037)) || ((pixel_index >= 3042) && (pixel_index <= 3099)) || ((pixel_index >= 3103) && (pixel_index <= 3134)) || ((pixel_index >= 3139) && (pixel_index <= 3195)) || ((pixel_index >= 3199) && (pixel_index <= 3231)) || ((pixel_index >= 3235) && (pixel_index <= 3291)) || ((pixel_index >= 3295) && (pixel_index <= 3327)) || ((pixel_index >= 3331) && (pixel_index <= 3387)) || ((pixel_index >= 3391) && (pixel_index <= 3424)) || ((pixel_index >= 3427) && (pixel_index <= 3483)) || ((pixel_index >= 3487) && (pixel_index <= 3520)) || ((pixel_index >= 3523) && (pixel_index <= 3580)) || ((pixel_index >= 3584) && (pixel_index <= 3616)) || ((pixel_index >= 3619) && (pixel_index <= 3676)) || ((pixel_index >= 3680) && (pixel_index <= 3712)) || ((pixel_index >= 3715) && (pixel_index <= 3773)) || ((pixel_index >= 3777) && (pixel_index <= 3807)) || ((pixel_index >= 3811) && (pixel_index <= 3869)) || ((pixel_index >= 3874) && (pixel_index <= 3885)) || ((pixel_index >= 3887) && (pixel_index <= 3903)) || ((pixel_index >= 3907) && (pixel_index <= 3966)) || ((pixel_index >= 3971) && (pixel_index <= 3979)) || ((pixel_index >= 3983) && (pixel_index <= 3986)) || ((pixel_index >= 3988) && (pixel_index <= 3998)) || ((pixel_index >= 4002) && (pixel_index <= 4063)) || ((pixel_index >= 4069) && (pixel_index <= 4073)) || ((pixel_index >= 4079) && (pixel_index <= 4082)) || ((pixel_index >= 4086) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4160)) || ((pixel_index >= 4174) && (pixel_index <= 4178)) || ((pixel_index >= 4192) && (pixel_index <= 4258)) || ((pixel_index >= 4267) && (pixel_index <= 4276)) || (pixel_index >= 4286) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2050 || pixel_index == 4173) oled_data = 16'b1010010100010100;
    else if (pixel_index == 3328) oled_data = 16'b1010011110010100;
    else oled_data = 0;
    end
    
    else if (freq>=554 && freq<587) //C#5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1389)) || ((pixel_index >= 1392) && (pixel_index <= 1395)) || ((pixel_index >= 1398) && (pixel_index <= 1485)) || ((pixel_index >= 1487) && (pixel_index <= 1491)) || ((pixel_index >= 1493) && (pixel_index <= 1581)) || ((pixel_index >= 1583) && (pixel_index <= 1587)) || ((pixel_index >= 1589) && (pixel_index <= 1676)) || ((pixel_index >= 1679) && (pixel_index <= 1682)) || ((pixel_index >= 1685) && (pixel_index <= 1755)) || ((pixel_index >= 1765) && (pixel_index <= 1772)) || ((pixel_index >= 1775) && (pixel_index <= 1778)) || ((pixel_index >= 1781) && (pixel_index <= 1786)) || ((pixel_index >= 1801) && (pixel_index <= 1849)) || ((pixel_index >= 1863) && (pixel_index <= 1866)) || ((pixel_index >= 1879) && (pixel_index <= 1882)) || ((pixel_index >= 1897) && (pixel_index <= 1944)) || ((pixel_index >= 1949) && (pixel_index <= 1955)) || ((pixel_index >= 1960) && (pixel_index <= 1964)) || ((pixel_index >= 1967) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 1978)) || ((pixel_index >= 1982) && (pixel_index <= 2039)) || ((pixel_index >= 2043) && (pixel_index <= 2053)) || ((pixel_index >= 2056) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2074)) || ((pixel_index >= 2078) && (pixel_index <= 2134)) || ((pixel_index >= 2138) && (pixel_index <= 2150)) || ((pixel_index >= 2152) && (pixel_index <= 2156)) || ((pixel_index >= 2159) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2170)) || ((pixel_index >= 2174) && (pixel_index <= 2230)) || ((pixel_index >= 2234) && (pixel_index <= 2252)) || ((pixel_index >= 2254) && (pixel_index <= 2258)) || ((pixel_index >= 2260) && (pixel_index <= 2266)) || ((pixel_index >= 2270) && (pixel_index <= 2325)) || ((pixel_index >= 2329) && (pixel_index <= 2348)) || ((pixel_index >= 2350) && (pixel_index <= 2354)) || ((pixel_index >= 2356) && (pixel_index <= 2362)) || ((pixel_index >= 2366) && (pixel_index <= 2421)) || ((pixel_index >= 2425) && (pixel_index <= 2441)) || ((pixel_index >= 2454) && (pixel_index <= 2458)) || ((pixel_index >= 2462) && (pixel_index <= 2516)) || ((pixel_index >= 2520) && (pixel_index <= 2537)) || ((pixel_index >= 2550) && (pixel_index <= 2554)) || ((pixel_index >= 2558) && (pixel_index <= 2612)) || ((pixel_index >= 2616) && (pixel_index <= 2635)) || ((pixel_index >= 2638) && (pixel_index <= 2641)) || ((pixel_index >= 2644) && (pixel_index <= 2650)) || ((pixel_index >= 2654) && (pixel_index <= 2708)) || ((pixel_index >= 2712) && (pixel_index <= 2731)) || ((pixel_index >= 2734) && (pixel_index <= 2737)) || ((pixel_index >= 2740) && (pixel_index <= 2746)) || ((pixel_index >= 2750) && (pixel_index <= 2804)) || ((pixel_index >= 2808) && (pixel_index <= 2827)) || ((pixel_index >= 2830) && (pixel_index <= 2833)) || ((pixel_index >= 2836) && (pixel_index <= 2842)) || ((pixel_index >= 2854) && (pixel_index <= 2900)) || ((pixel_index >= 2904) && (pixel_index <= 2923)) || ((pixel_index >= 2926) && (pixel_index <= 2929)) || ((pixel_index >= 2932) && (pixel_index <= 2939)) || ((pixel_index >= 2952) && (pixel_index <= 2996)) || ((pixel_index >= 3000) && (pixel_index <= 3019)) || ((pixel_index >= 3021) && (pixel_index <= 3025)) || ((pixel_index >= 3027) && (pixel_index <= 3044)) || ((pixel_index >= 3049) && (pixel_index <= 3092)) || ((pixel_index >= 3096) && (pixel_index <= 3141)) || ((pixel_index >= 3146) && (pixel_index <= 3188)) || ((pixel_index >= 3192) && (pixel_index <= 3238)) || ((pixel_index >= 3242) && (pixel_index <= 3284)) || ((pixel_index >= 3288) && (pixel_index <= 3335)) || ((pixel_index >= 3338) && (pixel_index <= 3380)) || ((pixel_index >= 3384) && (pixel_index <= 3431)) || ((pixel_index >= 3435) && (pixel_index <= 3476)) || ((pixel_index >= 3480) && (pixel_index <= 3527)) || ((pixel_index >= 3531) && (pixel_index <= 3573)) || ((pixel_index >= 3577) && (pixel_index <= 3623)) || ((pixel_index >= 3626) && (pixel_index <= 3669)) || ((pixel_index >= 3673) && (pixel_index <= 3719)) || ((pixel_index >= 3722) && (pixel_index <= 3765)) || ((pixel_index >= 3770) && (pixel_index <= 3814)) || ((pixel_index >= 3818) && (pixel_index <= 3862)) || ((pixel_index >= 3866) && (pixel_index <= 3878)) || ((pixel_index >= 3880) && (pixel_index <= 3910)) || ((pixel_index >= 3914) && (pixel_index <= 3959)) || ((pixel_index >= 3964) && (pixel_index <= 3972)) || ((pixel_index >= 3976) && (pixel_index <= 3993)) || ((pixel_index >= 3995) && (pixel_index <= 4005)) || ((pixel_index >= 4009) && (pixel_index <= 4056)) || ((pixel_index >= 4062) && (pixel_index <= 4066)) || ((pixel_index >= 4072) && (pixel_index <= 4089)) || ((pixel_index >= 4093) && (pixel_index <= 4099)) || ((pixel_index >= 4104) && (pixel_index <= 4153)) || ((pixel_index >= 4166) && (pixel_index <= 4185)) || ((pixel_index >= 4199) && (pixel_index <= 4251)) || ((pixel_index >= 4260) && (pixel_index <= 4283)) || (pixel_index >= 4293) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1397) oled_data = 16'b0000001010000000;
    else if (pixel_index == 1677 || pixel_index == 2164) oled_data = 16'b0101001010001010;
    else if (pixel_index == 1787 || pixel_index == 2931) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=587 && freq<622) //D5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1755)) || ((pixel_index >= 1768) && (pixel_index <= 1781)) || ((pixel_index >= 1795) && (pixel_index <= 1851)) || ((pixel_index >= 1866) && (pixel_index <= 1877)) || ((pixel_index >= 1891) && (pixel_index <= 1947)) || ((pixel_index >= 1951) && (pixel_index <= 1957)) || ((pixel_index >= 1964) && (pixel_index <= 1973)) || ((pixel_index >= 1976) && (pixel_index <= 2043)) || ((pixel_index >= 2047) && (pixel_index <= 2056)) || ((pixel_index >= 2061) && (pixel_index <= 2069)) || ((pixel_index >= 2072) && (pixel_index <= 2139)) || ((pixel_index >= 2143) && (pixel_index <= 2153)) || ((pixel_index >= 2158) && (pixel_index <= 2165)) || ((pixel_index >= 2168) && (pixel_index <= 2235)) || ((pixel_index >= 2239) && (pixel_index <= 2250)) || ((pixel_index >= 2254) && (pixel_index <= 2261)) || ((pixel_index >= 2264) && (pixel_index <= 2331)) || ((pixel_index >= 2335) && (pixel_index <= 2347)) || ((pixel_index >= 2351) && (pixel_index <= 2357)) || ((pixel_index >= 2360) && (pixel_index <= 2427)) || ((pixel_index >= 2431) && (pixel_index <= 2443)) || ((pixel_index >= 2447) && (pixel_index <= 2453)) || ((pixel_index >= 2456) && (pixel_index <= 2523)) || ((pixel_index >= 2527) && (pixel_index <= 2540)) || ((pixel_index >= 2543) && (pixel_index <= 2549)) || ((pixel_index >= 2552) && (pixel_index <= 2619)) || ((pixel_index >= 2623) && (pixel_index <= 2636)) || ((pixel_index >= 2640) && (pixel_index <= 2645)) || ((pixel_index >= 2648) && (pixel_index <= 2715)) || ((pixel_index >= 2719) && (pixel_index <= 2732)) || ((pixel_index >= 2736) && (pixel_index <= 2741)) || ((pixel_index >= 2744) && (pixel_index <= 2811)) || ((pixel_index >= 2815) && (pixel_index <= 2828)) || ((pixel_index >= 2832) && (pixel_index <= 2837)) || ((pixel_index >= 2849) && (pixel_index <= 2907)) || ((pixel_index >= 2911) && (pixel_index <= 2924)) || ((pixel_index >= 2928) && (pixel_index <= 2933)) || ((pixel_index >= 2946) && (pixel_index <= 3003)) || ((pixel_index >= 3007) && (pixel_index <= 3020)) || ((pixel_index >= 3024) && (pixel_index <= 3038)) || ((pixel_index >= 3043) && (pixel_index <= 3099)) || ((pixel_index >= 3103) && (pixel_index <= 3116)) || ((pixel_index >= 3120) && (pixel_index <= 3136)) || ((pixel_index >= 3140) && (pixel_index <= 3195)) || ((pixel_index >= 3199) && (pixel_index <= 3212)) || ((pixel_index >= 3216) && (pixel_index <= 3233)) || ((pixel_index >= 3237) && (pixel_index <= 3291)) || ((pixel_index >= 3295) && (pixel_index <= 3308)) || ((pixel_index >= 3312) && (pixel_index <= 3329)) || ((pixel_index >= 3333) && (pixel_index <= 3387)) || ((pixel_index >= 3391) && (pixel_index <= 3404)) || ((pixel_index >= 3408) && (pixel_index <= 3425)) || ((pixel_index >= 3429) && (pixel_index <= 3483)) || ((pixel_index >= 3487) && (pixel_index <= 3499)) || ((pixel_index >= 3503) && (pixel_index <= 3521)) || ((pixel_index >= 3525) && (pixel_index <= 3579)) || ((pixel_index >= 3583) && (pixel_index <= 3595)) || ((pixel_index >= 3599) && (pixel_index <= 3617)) || ((pixel_index >= 3621) && (pixel_index <= 3675)) || ((pixel_index >= 3679) && (pixel_index <= 3691)) || ((pixel_index >= 3695) && (pixel_index <= 3713)) || ((pixel_index >= 3717) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3786)) || ((pixel_index >= 3790) && (pixel_index <= 3809)) || ((pixel_index >= 3813) && (pixel_index <= 3867)) || ((pixel_index >= 3871) && (pixel_index <= 3881)) || ((pixel_index >= 3885) && (pixel_index <= 3904)) || ((pixel_index >= 3908) && (pixel_index <= 3963)) || ((pixel_index >= 3967) && (pixel_index <= 3975)) || ((pixel_index >= 3980) && (pixel_index <= 3987)) || ((pixel_index >= 3989) && (pixel_index <= 3999)) || ((pixel_index >= 4004) && (pixel_index <= 4059)) || ((pixel_index >= 4063) && (pixel_index <= 4067)) || ((pixel_index >= 4075) && (pixel_index <= 4083)) || ((pixel_index >= 4088) && (pixel_index <= 4093)) || ((pixel_index >= 4099) && (pixel_index <= 4155)) || ((pixel_index >= 4170) && (pixel_index <= 4180)) || ((pixel_index >= 4194) && (pixel_index <= 4251)) || ((pixel_index >= 4263) && (pixel_index <= 4278)) || (pixel_index >= 4288) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 3500 || pixel_index == 3812 || pixel_index == 4003 || pixel_index == 4068 || pixel_index == 4094 || pixel_index == 4193) oled_data = 16'b1010010100010100;
    else if (pixel_index == 4287) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=622 && freq<659) //Eb5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1290)) || ((pixel_index >= 1292) && (pixel_index <= 1386)) || ((pixel_index >= 1388) && (pixel_index <= 1482)) || ((pixel_index >= 1484) && (pixel_index <= 1578)) || ((pixel_index >= 1580) && (pixel_index <= 1674)) || ((pixel_index >= 1676) && (pixel_index <= 1750)) || ((pixel_index >= 1766) && (pixel_index <= 1770)) || ((pixel_index >= 1772) && (pixel_index <= 1786)) || ((pixel_index >= 1800) && (pixel_index <= 1846)) || ((pixel_index >= 1862) && (pixel_index <= 1866)) || ((pixel_index >= 1868) && (pixel_index <= 1869)) || ((pixel_index >= 1875) && (pixel_index <= 1882)) || ((pixel_index >= 1896) && (pixel_index <= 1942)) || ((pixel_index >= 1946) && (pixel_index <= 1962)) || pixel_index == 1964 || ((pixel_index >= 1967) && (pixel_index <= 1969)) || ((pixel_index >= 1972) && (pixel_index <= 1978)) || ((pixel_index >= 1981) && (pixel_index <= 2038)) || ((pixel_index >= 2042) && (pixel_index <= 2058)) || ((pixel_index >= 2061) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2074)) || ((pixel_index >= 2077) && (pixel_index <= 2134)) || ((pixel_index >= 2138) && (pixel_index <= 2154)) || ((pixel_index >= 2156) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2170)) || ((pixel_index >= 2173) && (pixel_index <= 2230)) || ((pixel_index >= 2234) && (pixel_index <= 2250)) || ((pixel_index >= 2252) && (pixel_index <= 2259)) || ((pixel_index >= 2261) && (pixel_index <= 2266)) || ((pixel_index >= 2269) && (pixel_index <= 2326)) || ((pixel_index >= 2330) && (pixel_index <= 2346)) || ((pixel_index >= 2348) && (pixel_index <= 2355)) || ((pixel_index >= 2358) && (pixel_index <= 2362)) || ((pixel_index >= 2365) && (pixel_index <= 2422)) || ((pixel_index >= 2426) && (pixel_index <= 2442)) || ((pixel_index >= 2444) && (pixel_index <= 2451)) || ((pixel_index >= 2454) && (pixel_index <= 2458)) || ((pixel_index >= 2461) && (pixel_index <= 2518)) || ((pixel_index >= 2522) && (pixel_index <= 2538)) || ((pixel_index >= 2540) && (pixel_index <= 2547)) || ((pixel_index >= 2549) && (pixel_index <= 2554)) || ((pixel_index >= 2557) && (pixel_index <= 2614)) || ((pixel_index >= 2618) && (pixel_index <= 2634)) || ((pixel_index >= 2636) && (pixel_index <= 2643)) || ((pixel_index >= 2645) && (pixel_index <= 2650)) || ((pixel_index >= 2653) && (pixel_index <= 2710)) || ((pixel_index >= 2714) && (pixel_index <= 2730)) || ((pixel_index >= 2732) && (pixel_index <= 2738)) || ((pixel_index >= 2741) && (pixel_index <= 2746)) || ((pixel_index >= 2749) && (pixel_index <= 2806)) || ((pixel_index >= 2810) && (pixel_index <= 2826)) || ((pixel_index >= 2829) && (pixel_index <= 2834)) || ((pixel_index >= 2837) && (pixel_index <= 2842)) || ((pixel_index >= 2854) && (pixel_index <= 2902)) || ((pixel_index >= 2916) && (pixel_index <= 2922)) || ((pixel_index >= 2927) && (pixel_index <= 2929)) || ((pixel_index >= 2932) && (pixel_index <= 2938)) || ((pixel_index >= 2951) && (pixel_index <= 2998)) || ((pixel_index >= 3012) && (pixel_index <= 3018)) || ((pixel_index >= 3020) && (pixel_index <= 3021)) || ((pixel_index >= 3027) && (pixel_index <= 3043)) || ((pixel_index >= 3048) && (pixel_index <= 3094)) || ((pixel_index >= 3098) && (pixel_index <= 3141)) || ((pixel_index >= 3145) && (pixel_index <= 3190)) || ((pixel_index >= 3194) && (pixel_index <= 3238)) || ((pixel_index >= 3241) && (pixel_index <= 3286)) || ((pixel_index >= 3290) && (pixel_index <= 3334)) || ((pixel_index >= 3338) && (pixel_index <= 3382)) || ((pixel_index >= 3386) && (pixel_index <= 3430)) || ((pixel_index >= 3434) && (pixel_index <= 3478)) || ((pixel_index >= 3482) && (pixel_index <= 3526)) || ((pixel_index >= 3530) && (pixel_index <= 3574)) || ((pixel_index >= 3578) && (pixel_index <= 3622)) || ((pixel_index >= 3626) && (pixel_index <= 3670)) || ((pixel_index >= 3674) && (pixel_index <= 3718)) || ((pixel_index >= 3722) && (pixel_index <= 3766)) || ((pixel_index >= 3770) && (pixel_index <= 3814)) || ((pixel_index >= 3817) && (pixel_index <= 3862)) || ((pixel_index >= 3866) && (pixel_index <= 3909)) || ((pixel_index >= 3913) && (pixel_index <= 3958)) || ((pixel_index >= 3962) && (pixel_index <= 3992)) || ((pixel_index >= 3994) && (pixel_index <= 4004)) || ((pixel_index >= 4008) && (pixel_index <= 4054)) || ((pixel_index >= 4058) && (pixel_index <= 4088)) || ((pixel_index >= 4093) && (pixel_index <= 4098)) || ((pixel_index >= 4104) && (pixel_index <= 4150)) || ((pixel_index >= 4166) && (pixel_index <= 4184)) || ((pixel_index >= 4198) && (pixel_index <= 4247)) || ((pixel_index >= 4262) && (pixel_index <= 4282)) || (pixel_index >= 4292) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1765 || pixel_index == 1861) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2357 || pixel_index == 4283) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=659 && freq<698) //E5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1758)) || ((pixel_index >= 1773) && (pixel_index <= 1778)) || ((pixel_index >= 1793) && (pixel_index <= 1854)) || ((pixel_index >= 1869) && (pixel_index <= 1874)) || ((pixel_index >= 1889) && (pixel_index <= 1950)) || ((pixel_index >= 1953) && (pixel_index <= 1970)) || ((pixel_index >= 1974) && (pixel_index <= 2046)) || ((pixel_index >= 2049) && (pixel_index <= 2066)) || ((pixel_index >= 2070) && (pixel_index <= 2142)) || ((pixel_index >= 2145) && (pixel_index <= 2162)) || ((pixel_index >= 2166) && (pixel_index <= 2238)) || ((pixel_index >= 2241) && (pixel_index <= 2258)) || ((pixel_index >= 2262) && (pixel_index <= 2334)) || ((pixel_index >= 2337) && (pixel_index <= 2354)) || ((pixel_index >= 2358) && (pixel_index <= 2430)) || ((pixel_index >= 2433) && (pixel_index <= 2450)) || ((pixel_index >= 2454) && (pixel_index <= 2526)) || ((pixel_index >= 2529) && (pixel_index <= 2546)) || ((pixel_index >= 2550) && (pixel_index <= 2622)) || ((pixel_index >= 2625) && (pixel_index <= 2642)) || ((pixel_index >= 2646) && (pixel_index <= 2718)) || ((pixel_index >= 2721) && (pixel_index <= 2738)) || ((pixel_index >= 2742) && (pixel_index <= 2814)) || ((pixel_index >= 2817) && (pixel_index <= 2834)) || ((pixel_index >= 2846) && (pixel_index <= 2910)) || ((pixel_index >= 2923) && (pixel_index <= 2930)) || ((pixel_index >= 2944) && (pixel_index <= 3006)) || ((pixel_index >= 3019) && (pixel_index <= 3036)) || ((pixel_index >= 3041) && (pixel_index <= 3102)) || ((pixel_index >= 3105) && (pixel_index <= 3133)) || ((pixel_index >= 3138) && (pixel_index <= 3198)) || ((pixel_index >= 3201) && (pixel_index <= 3230)) || ((pixel_index >= 3234) && (pixel_index <= 3294)) || ((pixel_index >= 3297) && (pixel_index <= 3327)) || ((pixel_index >= 3330) && (pixel_index <= 3390)) || ((pixel_index >= 3393) && (pixel_index <= 3423)) || ((pixel_index >= 3426) && (pixel_index <= 3486)) || ((pixel_index >= 3489) && (pixel_index <= 3519)) || ((pixel_index >= 3523) && (pixel_index <= 3582)) || ((pixel_index >= 3585) && (pixel_index <= 3615)) || ((pixel_index >= 3618) && (pixel_index <= 3678)) || ((pixel_index >= 3681) && (pixel_index <= 3711)) || ((pixel_index >= 3714) && (pixel_index <= 3774)) || ((pixel_index >= 3777) && (pixel_index <= 3806)) || ((pixel_index >= 3810) && (pixel_index <= 3870)) || ((pixel_index >= 3873) && (pixel_index <= 3902)) || ((pixel_index >= 3906) && (pixel_index <= 3966)) || ((pixel_index >= 3969) && (pixel_index <= 3985)) || ((pixel_index >= 3987) && (pixel_index <= 3997)) || ((pixel_index >= 4001) && (pixel_index <= 4062)) || ((pixel_index >= 4065) && (pixel_index <= 4081)) || ((pixel_index >= 4085) && (pixel_index <= 4091)) || ((pixel_index >= 4096) && (pixel_index <= 4158)) || ((pixel_index >= 4173) && (pixel_index <= 4177)) || ((pixel_index >= 4191) && (pixel_index <= 4254)) || ((pixel_index >= 4269) && (pixel_index <= 4275)) || (pixel_index >= 4285) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 3522) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=698 && freq<739) //F5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1758)) || ((pixel_index >= 1773) && (pixel_index <= 1778)) || ((pixel_index >= 1792) && (pixel_index <= 1854)) || ((pixel_index >= 1869) && (pixel_index <= 1874)) || ((pixel_index >= 1888) && (pixel_index <= 1950)) || ((pixel_index >= 1954) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 2046)) || ((pixel_index >= 2050) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2142)) || ((pixel_index >= 2146) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2238)) || ((pixel_index >= 2242) && (pixel_index <= 2258)) || ((pixel_index >= 2261) && (pixel_index <= 2334)) || ((pixel_index >= 2338) && (pixel_index <= 2354)) || ((pixel_index >= 2357) && (pixel_index <= 2430)) || ((pixel_index >= 2434) && (pixel_index <= 2450)) || ((pixel_index >= 2453) && (pixel_index <= 2526)) || ((pixel_index >= 2530) && (pixel_index <= 2546)) || ((pixel_index >= 2549) && (pixel_index <= 2622)) || ((pixel_index >= 2626) && (pixel_index <= 2642)) || ((pixel_index >= 2645) && (pixel_index <= 2718)) || ((pixel_index >= 2722) && (pixel_index <= 2738)) || ((pixel_index >= 2741) && (pixel_index <= 2814)) || ((pixel_index >= 2818) && (pixel_index <= 2834)) || ((pixel_index >= 2846) && (pixel_index <= 2910)) || ((pixel_index >= 2924) && (pixel_index <= 2930)) || ((pixel_index >= 2943) && (pixel_index <= 3006)) || ((pixel_index >= 3020) && (pixel_index <= 3035)) || ((pixel_index >= 3040) && (pixel_index <= 3102)) || ((pixel_index >= 3116) && (pixel_index <= 3133)) || ((pixel_index >= 3137) && (pixel_index <= 3198)) || ((pixel_index >= 3202) && (pixel_index <= 3229)) || ((pixel_index >= 3233) && (pixel_index <= 3294)) || ((pixel_index >= 3298) && (pixel_index <= 3326)) || ((pixel_index >= 3330) && (pixel_index <= 3390)) || ((pixel_index >= 3394) && (pixel_index <= 3422)) || ((pixel_index >= 3426) && (pixel_index <= 3486)) || ((pixel_index >= 3490) && (pixel_index <= 3518)) || ((pixel_index >= 3522) && (pixel_index <= 3582)) || ((pixel_index >= 3586) && (pixel_index <= 3614)) || ((pixel_index >= 3618) && (pixel_index <= 3678)) || ((pixel_index >= 3682) && (pixel_index <= 3710)) || ((pixel_index >= 3714) && (pixel_index <= 3774)) || ((pixel_index >= 3778) && (pixel_index <= 3806)) || ((pixel_index >= 3809) && (pixel_index <= 3870)) || ((pixel_index >= 3874) && (pixel_index <= 3901)) || ((pixel_index >= 3905) && (pixel_index <= 3966)) || ((pixel_index >= 3970) && (pixel_index <= 3984)) || ((pixel_index >= 3986) && (pixel_index <= 3996)) || ((pixel_index >= 4000) && (pixel_index <= 4062)) || ((pixel_index >= 4066) && (pixel_index <= 4080)) || ((pixel_index >= 4085) && (pixel_index <= 4090)) || ((pixel_index >= 4096) && (pixel_index <= 4158)) || ((pixel_index >= 4162) && (pixel_index <= 4176)) || ((pixel_index >= 4190) && (pixel_index <= 4254)) || ((pixel_index >= 4258) && (pixel_index <= 4274)) || (pixel_index >= 4284) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 3230 || pixel_index == 4275) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=739 && freq<784) //F#5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1387)) || ((pixel_index >= 1390) && (pixel_index <= 1393)) || ((pixel_index >= 1396) && (pixel_index <= 1483)) || ((pixel_index >= 1486) && (pixel_index <= 1489)) || ((pixel_index >= 1492) && (pixel_index <= 1579)) || ((pixel_index >= 1582) && (pixel_index <= 1585)) || ((pixel_index >= 1588) && (pixel_index <= 1675)) || ((pixel_index >= 1678) && (pixel_index <= 1681)) || ((pixel_index >= 1684) && (pixel_index <= 1751)) || ((pixel_index >= 1766) && (pixel_index <= 1771)) || ((pixel_index >= 1773) && (pixel_index <= 1777)) || ((pixel_index >= 1779) && (pixel_index <= 1785)) || ((pixel_index >= 1799) && (pixel_index <= 1847)) || ((pixel_index >= 1862) && (pixel_index <= 1864)) || ((pixel_index >= 1878) && (pixel_index <= 1881)) || ((pixel_index >= 1895) && (pixel_index <= 1943)) || ((pixel_index >= 1947) && (pixel_index <= 1962)) || ((pixel_index >= 1965) && (pixel_index <= 1968)) || ((pixel_index >= 1971) && (pixel_index <= 1977)) || ((pixel_index >= 1980) && (pixel_index <= 2039)) || ((pixel_index >= 2043) && (pixel_index <= 2058)) || ((pixel_index >= 2061) && (pixel_index <= 2064)) || ((pixel_index >= 2067) && (pixel_index <= 2073)) || ((pixel_index >= 2076) && (pixel_index <= 2135)) || ((pixel_index >= 2139) && (pixel_index <= 2154)) || ((pixel_index >= 2157) && (pixel_index <= 2160)) || ((pixel_index >= 2163) && (pixel_index <= 2169)) || ((pixel_index >= 2172) && (pixel_index <= 2231)) || ((pixel_index >= 2235) && (pixel_index <= 2250)) || ((pixel_index >= 2253) && (pixel_index <= 2256)) || ((pixel_index >= 2259) && (pixel_index <= 2265)) || ((pixel_index >= 2268) && (pixel_index <= 2327)) || ((pixel_index >= 2331) && (pixel_index <= 2346)) || ((pixel_index >= 2349) && (pixel_index <= 2352)) || ((pixel_index >= 2355) && (pixel_index <= 2361)) || ((pixel_index >= 2364) && (pixel_index <= 2423)) || ((pixel_index >= 2427) && (pixel_index <= 2440)) || ((pixel_index >= 2453) && (pixel_index <= 2457)) || ((pixel_index >= 2460) && (pixel_index <= 2519)) || ((pixel_index >= 2523) && (pixel_index <= 2535)) || ((pixel_index >= 2549) && (pixel_index <= 2553)) || ((pixel_index >= 2556) && (pixel_index <= 2615)) || ((pixel_index >= 2619) && (pixel_index <= 2634)) || ((pixel_index >= 2636) && (pixel_index <= 2640)) || ((pixel_index >= 2642) && (pixel_index <= 2649)) || ((pixel_index >= 2652) && (pixel_index <= 2711)) || ((pixel_index >= 2715) && (pixel_index <= 2729)) || ((pixel_index >= 2732) && (pixel_index <= 2735)) || ((pixel_index >= 2738) && (pixel_index <= 2745)) || ((pixel_index >= 2748) && (pixel_index <= 2807)) || ((pixel_index >= 2811) && (pixel_index <= 2825)) || ((pixel_index >= 2828) && (pixel_index <= 2831)) || ((pixel_index >= 2834) && (pixel_index <= 2841)) || ((pixel_index >= 2853) && (pixel_index <= 2903)) || ((pixel_index >= 2917) && (pixel_index <= 2921)) || ((pixel_index >= 2924) && (pixel_index <= 2927)) || ((pixel_index >= 2930) && (pixel_index <= 2937)) || ((pixel_index >= 2950) && (pixel_index <= 2999)) || ((pixel_index >= 3013) && (pixel_index <= 3017)) || ((pixel_index >= 3020) && (pixel_index <= 3023)) || ((pixel_index >= 3026) && (pixel_index <= 3042)) || ((pixel_index >= 3047) && (pixel_index <= 3095)) || ((pixel_index >= 3109) && (pixel_index <= 3140)) || ((pixel_index >= 3144) && (pixel_index <= 3191)) || ((pixel_index >= 3195) && (pixel_index <= 3237)) || ((pixel_index >= 3241) && (pixel_index <= 3287)) || ((pixel_index >= 3291) && (pixel_index <= 3333)) || ((pixel_index >= 3337) && (pixel_index <= 3383)) || ((pixel_index >= 3387) && (pixel_index <= 3429)) || ((pixel_index >= 3433) && (pixel_index <= 3479)) || ((pixel_index >= 3483) && (pixel_index <= 3525)) || ((pixel_index >= 3529) && (pixel_index <= 3575)) || ((pixel_index >= 3579) && (pixel_index <= 3621)) || ((pixel_index >= 3625) && (pixel_index <= 3671)) || ((pixel_index >= 3675) && (pixel_index <= 3717)) || ((pixel_index >= 3721) && (pixel_index <= 3767)) || ((pixel_index >= 3771) && (pixel_index <= 3813)) || ((pixel_index >= 3816) && (pixel_index <= 3863)) || ((pixel_index >= 3867) && (pixel_index <= 3908)) || ((pixel_index >= 3912) && (pixel_index <= 3959)) || ((pixel_index >= 3963) && (pixel_index <= 3991)) || ((pixel_index >= 3993) && (pixel_index <= 4003)) || ((pixel_index >= 4007) && (pixel_index <= 4055)) || ((pixel_index >= 4059) && (pixel_index <= 4087)) || ((pixel_index >= 4092) && (pixel_index <= 4097)) || ((pixel_index >= 4103) && (pixel_index <= 4151)) || ((pixel_index >= 4155) && (pixel_index <= 4183)) || ((pixel_index >= 4197) && (pixel_index <= 4247)) || ((pixel_index >= 4251) && (pixel_index <= 4281)) || (pixel_index >= 4292) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1963 || pixel_index == 3240 || pixel_index == 4184) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2536) oled_data = 16'b1010011110010100;
    else if (pixel_index == 4282 || pixel_index == 4291) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=784 && freq<830) //G5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1761)) || ((pixel_index >= 1772) && (pixel_index <= 1781)) || ((pixel_index >= 1796) && (pixel_index <= 1855)) || ((pixel_index >= 1870) && (pixel_index <= 1877)) || ((pixel_index >= 1892) && (pixel_index <= 1949)) || ((pixel_index >= 1955) && (pixel_index <= 1962)) || ((pixel_index >= 1967) && (pixel_index <= 1973)) || ((pixel_index >= 1977) && (pixel_index <= 2044)) || ((pixel_index >= 2049) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2069)) || ((pixel_index >= 2073) && (pixel_index <= 2140)) || ((pixel_index >= 2144) && (pixel_index <= 2165)) || ((pixel_index >= 2169) && (pixel_index <= 2235)) || ((pixel_index >= 2239) && (pixel_index <= 2261)) || ((pixel_index >= 2265) && (pixel_index <= 2330)) || ((pixel_index >= 2334) && (pixel_index <= 2357)) || ((pixel_index >= 2361) && (pixel_index <= 2426)) || ((pixel_index >= 2430) && (pixel_index <= 2453)) || ((pixel_index >= 2457) && (pixel_index <= 2522)) || ((pixel_index >= 2525) && (pixel_index <= 2549)) || ((pixel_index >= 2553) && (pixel_index <= 2617)) || ((pixel_index >= 2621) && (pixel_index <= 2645)) || ((pixel_index >= 2649) && (pixel_index <= 2713)) || ((pixel_index >= 2717) && (pixel_index <= 2741)) || ((pixel_index >= 2745) && (pixel_index <= 2809)) || ((pixel_index >= 2813) && (pixel_index <= 2837)) || ((pixel_index >= 2849) && (pixel_index <= 2905)) || ((pixel_index >= 2909) && (pixel_index <= 2916)) || ((pixel_index >= 2927) && (pixel_index <= 2933)) || ((pixel_index >= 2947) && (pixel_index <= 3001)) || ((pixel_index >= 3005) && (pixel_index <= 3012)) || ((pixel_index >= 3023) && (pixel_index <= 3039)) || ((pixel_index >= 3044) && (pixel_index <= 3097)) || ((pixel_index >= 3101) && (pixel_index <= 3108)) || ((pixel_index >= 3119) && (pixel_index <= 3136)) || ((pixel_index >= 3141) && (pixel_index <= 3193)) || ((pixel_index >= 3197) && (pixel_index <= 3212)) || ((pixel_index >= 3215) && (pixel_index <= 3233)) || ((pixel_index >= 3237) && (pixel_index <= 3289)) || ((pixel_index >= 3293) && (pixel_index <= 3308)) || ((pixel_index >= 3311) && (pixel_index <= 3329)) || ((pixel_index >= 3333) && (pixel_index <= 3385)) || ((pixel_index >= 3389) && (pixel_index <= 3404)) || ((pixel_index >= 3407) && (pixel_index <= 3426)) || ((pixel_index >= 3429) && (pixel_index <= 3482)) || ((pixel_index >= 3486) && (pixel_index <= 3500)) || ((pixel_index >= 3503) && (pixel_index <= 3522)) || ((pixel_index >= 3525) && (pixel_index <= 3578)) || ((pixel_index >= 3582) && (pixel_index <= 3596)) || ((pixel_index >= 3599) && (pixel_index <= 3618)) || ((pixel_index >= 3621) && (pixel_index <= 3674)) || ((pixel_index >= 3679) && (pixel_index <= 3692)) || ((pixel_index >= 3695) && (pixel_index <= 3714)) || ((pixel_index >= 3717) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3788)) || ((pixel_index >= 3791) && (pixel_index <= 3809)) || ((pixel_index >= 3813) && (pixel_index <= 3868)) || ((pixel_index >= 3872) && (pixel_index <= 3884)) || ((pixel_index >= 3887) && (pixel_index <= 3905)) || ((pixel_index >= 3909) && (pixel_index <= 3964)) || ((pixel_index >= 3970) && (pixel_index <= 3979)) || ((pixel_index >= 3983) && (pixel_index <= 3988)) || ((pixel_index >= 3990) && (pixel_index <= 4000)) || ((pixel_index >= 4004) && (pixel_index <= 4061)) || ((pixel_index >= 4068) && (pixel_index <= 4073)) || ((pixel_index >= 4079) && (pixel_index <= 4084)) || ((pixel_index >= 4088) && (pixel_index <= 4094)) || ((pixel_index >= 4099) && (pixel_index <= 4159)) || ((pixel_index >= 4174) && (pixel_index <= 4180)) || ((pixel_index >= 4194) && (pixel_index <= 4257)) || ((pixel_index >= 4267) && (pixel_index <= 4278)) || (pixel_index >= 4288) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2926 || pixel_index == 3330 || pixel_index == 3485 || pixel_index == 3678) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=830 && freq<880) //Ab5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1291)) || ((pixel_index >= 1294) && (pixel_index <= 1387)) || ((pixel_index >= 1390) && (pixel_index <= 1483)) || ((pixel_index >= 1486) && (pixel_index <= 1579)) || ((pixel_index >= 1582) && (pixel_index <= 1675)) || ((pixel_index >= 1678) && (pixel_index <= 1755)) || ((pixel_index >= 1759) && (pixel_index <= 1771)) || ((pixel_index >= 1774) && (pixel_index <= 1787)) || ((pixel_index >= 1802) && (pixel_index <= 1851)) || ((pixel_index >= 1856) && (pixel_index <= 1867)) || pixel_index == 1870 || ((pixel_index >= 1877) && (pixel_index <= 1883)) || ((pixel_index >= 1898) && (pixel_index <= 1946)) || ((pixel_index >= 1952) && (pixel_index <= 1963)) || ((pixel_index >= 1968) && (pixel_index <= 1970)) || ((pixel_index >= 1974) && (pixel_index <= 1979)) || ((pixel_index >= 1983) && (pixel_index <= 2042)) || pixel_index == 2045 || ((pixel_index >= 2049) && (pixel_index <= 2059)) || ((pixel_index >= 2063) && (pixel_index <= 2067)) || ((pixel_index >= 2070) && (pixel_index <= 2075)) || ((pixel_index >= 2079) && (pixel_index <= 2138)) || pixel_index == 2141 || ((pixel_index >= 2145) && (pixel_index <= 2155)) || ((pixel_index >= 2158) && (pixel_index <= 2164)) || ((pixel_index >= 2167) && (pixel_index <= 2171)) || ((pixel_index >= 2175) && (pixel_index <= 2233)) || ((pixel_index >= 2237) && (pixel_index <= 2238)) || ((pixel_index >= 2241) && (pixel_index <= 2251)) || ((pixel_index >= 2254) && (pixel_index <= 2260)) || ((pixel_index >= 2263) && (pixel_index <= 2267)) || ((pixel_index >= 2271) && (pixel_index <= 2329)) || ((pixel_index >= 2332) && (pixel_index <= 2334)) || ((pixel_index >= 2338) && (pixel_index <= 2347)) || ((pixel_index >= 2350) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2363)) || ((pixel_index >= 2367) && (pixel_index <= 2424)) || ((pixel_index >= 2428) && (pixel_index <= 2430)) || ((pixel_index >= 2434) && (pixel_index <= 2443)) || ((pixel_index >= 2446) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2459)) || ((pixel_index >= 2463) && (pixel_index <= 2520)) || ((pixel_index >= 2524) && (pixel_index <= 2527)) || ((pixel_index >= 2530) && (pixel_index <= 2539)) || ((pixel_index >= 2542) && (pixel_index <= 2548)) || ((pixel_index >= 2551) && (pixel_index <= 2555)) || ((pixel_index >= 2559) && (pixel_index <= 2616)) || ((pixel_index >= 2619) && (pixel_index <= 2623)) || ((pixel_index >= 2627) && (pixel_index <= 2635)) || ((pixel_index >= 2638) && (pixel_index <= 2644)) || ((pixel_index >= 2647) && (pixel_index <= 2651)) || ((pixel_index >= 2655) && (pixel_index <= 2711)) || ((pixel_index >= 2715) && (pixel_index <= 2719)) || ((pixel_index >= 2723) && (pixel_index <= 2731)) || ((pixel_index >= 2734) && (pixel_index <= 2740)) || ((pixel_index >= 2743) && (pixel_index <= 2747)) || ((pixel_index >= 2751) && (pixel_index <= 2807)) || ((pixel_index >= 2810) && (pixel_index <= 2816)) || ((pixel_index >= 2820) && (pixel_index <= 2827)) || ((pixel_index >= 2831) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2843)) || ((pixel_index >= 2855) && (pixel_index <= 2903)) || ((pixel_index >= 2906) && (pixel_index <= 2912)) || ((pixel_index >= 2916) && (pixel_index <= 2923)) || ((pixel_index >= 2928) && (pixel_index <= 2930)) || ((pixel_index >= 2934) && (pixel_index <= 2939)) || ((pixel_index >= 2953) && (pixel_index <= 2998)) || ((pixel_index >= 3002) && (pixel_index <= 3009)) || ((pixel_index >= 3012) && (pixel_index <= 3019)) || pixel_index == 3022 || ((pixel_index >= 3029) && (pixel_index <= 3045)) || ((pixel_index >= 3050) && (pixel_index <= 3094)) || ((pixel_index >= 3097) && (pixel_index <= 3105)) || ((pixel_index >= 3109) && (pixel_index <= 3142)) || ((pixel_index >= 3147) && (pixel_index <= 3190)) || ((pixel_index >= 3193) && (pixel_index <= 3201)) || ((pixel_index >= 3205) && (pixel_index <= 3239)) || ((pixel_index >= 3243) && (pixel_index <= 3285)) || ((pixel_index >= 3289) && (pixel_index <= 3298)) || ((pixel_index >= 3301) && (pixel_index <= 3336)) || ((pixel_index >= 3339) && (pixel_index <= 3381)) || ((pixel_index >= 3398) && (pixel_index <= 3432)) || ((pixel_index >= 3435) && (pixel_index <= 3476)) || ((pixel_index >= 3494) && (pixel_index <= 3528)) || ((pixel_index >= 3531) && (pixel_index <= 3572)) || ((pixel_index >= 3576) && (pixel_index <= 3587)) || ((pixel_index >= 3590) && (pixel_index <= 3624)) || ((pixel_index >= 3627) && (pixel_index <= 3668)) || ((pixel_index >= 3671) && (pixel_index <= 3683)) || ((pixel_index >= 3687) && (pixel_index <= 3720)) || ((pixel_index >= 3723) && (pixel_index <= 3763)) || ((pixel_index >= 3767) && (pixel_index <= 3779)) || ((pixel_index >= 3783) && (pixel_index <= 3815)) || ((pixel_index >= 3819) && (pixel_index <= 3859)) || ((pixel_index >= 3863) && (pixel_index <= 3876)) || ((pixel_index >= 3880) && (pixel_index <= 3911)) || ((pixel_index >= 3915) && (pixel_index <= 3955)) || ((pixel_index >= 3958) && (pixel_index <= 3972)) || ((pixel_index >= 3976) && (pixel_index <= 3994)) || ((pixel_index >= 3996) && (pixel_index <= 4006)) || ((pixel_index >= 4010) && (pixel_index <= 4050)) || ((pixel_index >= 4054) && (pixel_index <= 4068)) || ((pixel_index >= 4072) && (pixel_index <= 4090)) || ((pixel_index >= 4094) && (pixel_index <= 4100)) || ((pixel_index >= 4105) && (pixel_index <= 4146)) || ((pixel_index >= 4150) && (pixel_index <= 4165)) || ((pixel_index >= 4169) && (pixel_index <= 4186)) || ((pixel_index >= 4200) && (pixel_index <= 4242)) || ((pixel_index >= 4245) && (pixel_index <= 4261)) || ((pixel_index >= 4265) && (pixel_index <= 4284)) || (pixel_index >= 4294) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1971) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2819) oled_data = 16'b0101010100001010;
    else if (pixel_index == 4069) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=880 && freq<932) //A5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1762)) || ((pixel_index >= 1767) && (pixel_index <= 1780)) || ((pixel_index >= 1794) && (pixel_index <= 1858)) || ((pixel_index >= 1863) && (pixel_index <= 1876)) || ((pixel_index >= 1890) && (pixel_index <= 1954)) || ((pixel_index >= 1960) && (pixel_index <= 1972)) || ((pixel_index >= 1975) && (pixel_index <= 2049)) || ((pixel_index >= 2056) && (pixel_index <= 2068)) || ((pixel_index >= 2071) && (pixel_index <= 2145)) || ((pixel_index >= 2148) && (pixel_index <= 2149)) || ((pixel_index >= 2152) && (pixel_index <= 2164)) || ((pixel_index >= 2167) && (pixel_index <= 2241)) || ((pixel_index >= 2244) && (pixel_index <= 2245)) || ((pixel_index >= 2249) && (pixel_index <= 2260)) || ((pixel_index >= 2263) && (pixel_index <= 2336)) || ((pixel_index >= 2340) && (pixel_index <= 2341)) || ((pixel_index >= 2345) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2432)) || ((pixel_index >= 2435) && (pixel_index <= 2438)) || ((pixel_index >= 2441) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2527)) || ((pixel_index >= 2531) && (pixel_index <= 2534)) || ((pixel_index >= 2538) && (pixel_index <= 2548)) || ((pixel_index >= 2551) && (pixel_index <= 2623)) || ((pixel_index >= 2627) && (pixel_index <= 2630)) || ((pixel_index >= 2634) && (pixel_index <= 2644)) || ((pixel_index >= 2647) && (pixel_index <= 2719)) || ((pixel_index >= 2722) && (pixel_index <= 2727)) || ((pixel_index >= 2731) && (pixel_index <= 2740)) || ((pixel_index >= 2743) && (pixel_index <= 2814)) || ((pixel_index >= 2818) && (pixel_index <= 2823)) || ((pixel_index >= 2827) && (pixel_index <= 2836)) || ((pixel_index >= 2848) && (pixel_index <= 2910)) || ((pixel_index >= 2914) && (pixel_index <= 2920)) || ((pixel_index >= 2923) && (pixel_index <= 2932)) || ((pixel_index >= 2946) && (pixel_index <= 3006)) || ((pixel_index >= 3009) && (pixel_index <= 3016)) || ((pixel_index >= 3020) && (pixel_index <= 3037)) || ((pixel_index >= 3043) && (pixel_index <= 3101)) || ((pixel_index >= 3105) && (pixel_index <= 3112)) || ((pixel_index >= 3116) && (pixel_index <= 3135)) || ((pixel_index >= 3139) && (pixel_index <= 3197)) || ((pixel_index >= 3201) && (pixel_index <= 3209)) || ((pixel_index >= 3212) && (pixel_index <= 3232)) || ((pixel_index >= 3236) && (pixel_index <= 3293)) || ((pixel_index >= 3296) && (pixel_index <= 3305)) || ((pixel_index >= 3309) && (pixel_index <= 3328)) || ((pixel_index >= 3332) && (pixel_index <= 3388)) || ((pixel_index >= 3405) && (pixel_index <= 3424)) || ((pixel_index >= 3428) && (pixel_index <= 3484)) || ((pixel_index >= 3501) && (pixel_index <= 3520)) || ((pixel_index >= 3524) && (pixel_index <= 3579)) || ((pixel_index >= 3583) && (pixel_index <= 3594)) || ((pixel_index >= 3598) && (pixel_index <= 3616)) || ((pixel_index >= 3620) && (pixel_index <= 3675)) || ((pixel_index >= 3679) && (pixel_index <= 3690)) || ((pixel_index >= 3694) && (pixel_index <= 3712)) || ((pixel_index >= 3716) && (pixel_index <= 3771)) || ((pixel_index >= 3774) && (pixel_index <= 3787)) || ((pixel_index >= 3791) && (pixel_index <= 3808)) || ((pixel_index >= 3812) && (pixel_index <= 3866)) || ((pixel_index >= 3870) && (pixel_index <= 3883)) || ((pixel_index >= 3887) && (pixel_index <= 3903)) || ((pixel_index >= 3907) && (pixel_index <= 3962)) || ((pixel_index >= 3966) && (pixel_index <= 3980)) || ((pixel_index >= 3983) && (pixel_index <= 3987)) || ((pixel_index >= 3989) && (pixel_index <= 3998)) || ((pixel_index >= 4003) && (pixel_index <= 4058)) || ((pixel_index >= 4061) && (pixel_index <= 4076)) || ((pixel_index >= 4080) && (pixel_index <= 4082)) || ((pixel_index >= 4087) && (pixel_index <= 4093)) || ((pixel_index >= 4098) && (pixel_index <= 4153)) || ((pixel_index >= 4157) && (pixel_index <= 4172)) || ((pixel_index >= 4176) && (pixel_index <= 4179)) || ((pixel_index >= 4193) && (pixel_index <= 4249)) || ((pixel_index >= 4253) && (pixel_index <= 4269)) || ((pixel_index >= 4272) && (pixel_index <= 4277)) || (pixel_index >= 4287) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2528 || pixel_index == 2631 || pixel_index == 3200) oled_data = 16'b1010010100010100;
    else if (pixel_index == 3038) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=932 && freq<987) //Bb5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1290)) || ((pixel_index >= 1293) && (pixel_index <= 1386)) || ((pixel_index >= 1389) && (pixel_index <= 1482)) || ((pixel_index >= 1485) && (pixel_index <= 1578)) || ((pixel_index >= 1581) && (pixel_index <= 1674)) || ((pixel_index >= 1677) && (pixel_index <= 1749)) || ((pixel_index >= 1762) && (pixel_index <= 1770)) || ((pixel_index >= 1773) && (pixel_index <= 1787)) || ((pixel_index >= 1801) && (pixel_index <= 1845)) || ((pixel_index >= 1859) && (pixel_index <= 1866)) || ((pixel_index >= 1869) && (pixel_index <= 1870)) || ((pixel_index >= 1876) && (pixel_index <= 1883)) || ((pixel_index >= 1897) && (pixel_index <= 1941)) || ((pixel_index >= 1945) && (pixel_index <= 1951)) || ((pixel_index >= 1956) && (pixel_index <= 1962)) || ((pixel_index >= 1968) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 1979)) || ((pixel_index >= 1982) && (pixel_index <= 2037)) || ((pixel_index >= 2041) && (pixel_index <= 2048)) || ((pixel_index >= 2053) && (pixel_index <= 2058)) || ((pixel_index >= 2062) && (pixel_index <= 2067)) || ((pixel_index >= 2070) && (pixel_index <= 2075)) || ((pixel_index >= 2078) && (pixel_index <= 2133)) || ((pixel_index >= 2137) && (pixel_index <= 2145)) || ((pixel_index >= 2149) && (pixel_index <= 2154)) || ((pixel_index >= 2157) && (pixel_index <= 2163)) || ((pixel_index >= 2166) && (pixel_index <= 2171)) || ((pixel_index >= 2174) && (pixel_index <= 2229)) || ((pixel_index >= 2233) && (pixel_index <= 2241)) || ((pixel_index >= 2245) && (pixel_index <= 2250)) || ((pixel_index >= 2253) && (pixel_index <= 2260)) || ((pixel_index >= 2262) && (pixel_index <= 2267)) || ((pixel_index >= 2270) && (pixel_index <= 2325)) || ((pixel_index >= 2329) && (pixel_index <= 2338)) || ((pixel_index >= 2341) && (pixel_index <= 2346)) || ((pixel_index >= 2349) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2363)) || ((pixel_index >= 2366) && (pixel_index <= 2421)) || ((pixel_index >= 2425) && (pixel_index <= 2434)) || ((pixel_index >= 2437) && (pixel_index <= 2442)) || ((pixel_index >= 2445) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2459)) || ((pixel_index >= 2462) && (pixel_index <= 2517)) || ((pixel_index >= 2521) && (pixel_index <= 2529)) || ((pixel_index >= 2533) && (pixel_index <= 2538)) || ((pixel_index >= 2541) && (pixel_index <= 2548)) || ((pixel_index >= 2550) && (pixel_index <= 2555)) || ((pixel_index >= 2558) && (pixel_index <= 2613)) || ((pixel_index >= 2617) && (pixel_index <= 2625)) || ((pixel_index >= 2629) && (pixel_index <= 2634)) || ((pixel_index >= 2637) && (pixel_index <= 2644)) || ((pixel_index >= 2646) && (pixel_index <= 2651)) || ((pixel_index >= 2654) && (pixel_index <= 2709)) || ((pixel_index >= 2713) && (pixel_index <= 2720)) || ((pixel_index >= 2724) && (pixel_index <= 2730)) || ((pixel_index >= 2733) && (pixel_index <= 2739)) || ((pixel_index >= 2742) && (pixel_index <= 2747)) || ((pixel_index >= 2750) && (pixel_index <= 2805)) || ((pixel_index >= 2809) && (pixel_index <= 2815)) || ((pixel_index >= 2819) && (pixel_index <= 2826)) || ((pixel_index >= 2830) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2843)) || ((pixel_index >= 2855) && (pixel_index <= 2901)) || ((pixel_index >= 2914) && (pixel_index <= 2922)) || ((pixel_index >= 2928) && (pixel_index <= 2930)) || ((pixel_index >= 2933) && (pixel_index <= 2939)) || ((pixel_index >= 2952) && (pixel_index <= 2997)) || ((pixel_index >= 3012) && (pixel_index <= 3018)) || ((pixel_index >= 3021) && (pixel_index <= 3022)) || ((pixel_index >= 3028) && (pixel_index <= 3044)) || ((pixel_index >= 3049) && (pixel_index <= 3093)) || ((pixel_index >= 3097) && (pixel_index <= 3104)) || ((pixel_index >= 3109) && (pixel_index <= 3142)) || ((pixel_index >= 3146) && (pixel_index <= 3189)) || ((pixel_index >= 3193) && (pixel_index <= 3202)) || ((pixel_index >= 3206) && (pixel_index <= 3238)) || ((pixel_index >= 3242) && (pixel_index <= 3285)) || ((pixel_index >= 3289) && (pixel_index <= 3299)) || ((pixel_index >= 3303) && (pixel_index <= 3335)) || ((pixel_index >= 3339) && (pixel_index <= 3381)) || ((pixel_index >= 3385) && (pixel_index <= 3395)) || ((pixel_index >= 3399) && (pixel_index <= 3431)) || ((pixel_index >= 3435) && (pixel_index <= 3477)) || ((pixel_index >= 3481) && (pixel_index <= 3491)) || ((pixel_index >= 3495) && (pixel_index <= 3527)) || ((pixel_index >= 3531) && (pixel_index <= 3573)) || ((pixel_index >= 3577) && (pixel_index <= 3587)) || ((pixel_index >= 3591) && (pixel_index <= 3623)) || ((pixel_index >= 3627) && (pixel_index <= 3669)) || ((pixel_index >= 3673) && (pixel_index <= 3683)) || ((pixel_index >= 3687) && (pixel_index <= 3719)) || ((pixel_index >= 3723) && (pixel_index <= 3765)) || ((pixel_index >= 3769) && (pixel_index <= 3779)) || ((pixel_index >= 3783) && (pixel_index <= 3815)) || ((pixel_index >= 3818) && (pixel_index <= 3861)) || ((pixel_index >= 3865) && (pixel_index <= 3874)) || ((pixel_index >= 3878) && (pixel_index <= 3910)) || ((pixel_index >= 3914) && (pixel_index <= 3957)) || ((pixel_index >= 3961) && (pixel_index <= 3969)) || ((pixel_index >= 3974) && (pixel_index <= 3993)) || ((pixel_index >= 3995) && (pixel_index <= 4005)) || ((pixel_index >= 4009) && (pixel_index <= 4053)) || ((pixel_index >= 4057) && (pixel_index <= 4063)) || ((pixel_index >= 4069) && (pixel_index <= 4089)) || ((pixel_index >= 4094) && (pixel_index <= 4099)) || ((pixel_index >= 4105) && (pixel_index <= 4149)) || ((pixel_index >= 4164) && (pixel_index <= 4185)) || ((pixel_index >= 4199) && (pixel_index <= 4246)) || ((pixel_index >= 4258) && (pixel_index <= 4283)) || (pixel_index >= 4293) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1291 || pixel_index == 1387 || pixel_index == 1483 || pixel_index == 1579 || pixel_index == 1675 || pixel_index == 1771 || pixel_index == 1867 || pixel_index == 1963 || pixel_index == 1965 || pixel_index == 2059 || pixel_index == 2155 || pixel_index == 2251 || pixel_index == 2347 || pixel_index == 2358 || pixel_index == 2443 || pixel_index == 2539 || pixel_index == 2635 || pixel_index == 2731 || pixel_index == 2827 || pixel_index == 2923 || pixel_index == 3019 || pixel_index == 3239) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2049 || pixel_index == 2242 || pixel_index == 4284) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=987 && freq<1046) //B5
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1757)) || ((pixel_index >= 1769) && (pixel_index <= 1779)) || ((pixel_index >= 1794) && (pixel_index <= 1853)) || ((pixel_index >= 1867) && (pixel_index <= 1875)) || ((pixel_index >= 1890) && (pixel_index <= 1949)) || ((pixel_index >= 1952) && (pixel_index <= 1958)) || ((pixel_index >= 1964) && (pixel_index <= 1971)) || ((pixel_index >= 1975) && (pixel_index <= 2045)) || ((pixel_index >= 2048) && (pixel_index <= 2056)) || ((pixel_index >= 2060) && (pixel_index <= 2067)) || ((pixel_index >= 2071) && (pixel_index <= 2141)) || ((pixel_index >= 2144) && (pixel_index <= 2153)) || ((pixel_index >= 2157) && (pixel_index <= 2163)) || ((pixel_index >= 2167) && (pixel_index <= 2237)) || ((pixel_index >= 2240) && (pixel_index <= 2249)) || ((pixel_index >= 2253) && (pixel_index <= 2259)) || ((pixel_index >= 2263) && (pixel_index <= 2333)) || ((pixel_index >= 2336) && (pixel_index <= 2345)) || ((pixel_index >= 2349) && (pixel_index <= 2355)) || ((pixel_index >= 2359) && (pixel_index <= 2429)) || ((pixel_index >= 2432) && (pixel_index <= 2441)) || ((pixel_index >= 2445) && (pixel_index <= 2451)) || ((pixel_index >= 2455) && (pixel_index <= 2525)) || ((pixel_index >= 2528) && (pixel_index <= 2537)) || ((pixel_index >= 2541) && (pixel_index <= 2547)) || ((pixel_index >= 2551) && (pixel_index <= 2621)) || ((pixel_index >= 2624) && (pixel_index <= 2632)) || ((pixel_index >= 2636) && (pixel_index <= 2643)) || ((pixel_index >= 2647) && (pixel_index <= 2717)) || ((pixel_index >= 2720) && (pixel_index <= 2728)) || ((pixel_index >= 2732) && (pixel_index <= 2739)) || ((pixel_index >= 2743) && (pixel_index <= 2813)) || ((pixel_index >= 2816) && (pixel_index <= 2822)) || ((pixel_index >= 2827) && (pixel_index <= 2835)) || ((pixel_index >= 2847) && (pixel_index <= 2909)) || ((pixel_index >= 2921) && (pixel_index <= 2931)) || ((pixel_index >= 2945) && (pixel_index <= 3005)) || ((pixel_index >= 3020) && (pixel_index <= 3037)) || ((pixel_index >= 3042) && (pixel_index <= 3101)) || ((pixel_index >= 3104) && (pixel_index <= 3111)) || ((pixel_index >= 3117) && (pixel_index <= 3134)) || ((pixel_index >= 3139) && (pixel_index <= 3197)) || ((pixel_index >= 3200) && (pixel_index <= 3209)) || ((pixel_index >= 3214) && (pixel_index <= 3231)) || ((pixel_index >= 3235) && (pixel_index <= 3293)) || ((pixel_index >= 3296) && (pixel_index <= 3306)) || ((pixel_index >= 3310) && (pixel_index <= 3327)) || ((pixel_index >= 3331) && (pixel_index <= 3389)) || ((pixel_index >= 3392) && (pixel_index <= 3402)) || ((pixel_index >= 3406) && (pixel_index <= 3424)) || ((pixel_index >= 3427) && (pixel_index <= 3485)) || ((pixel_index >= 3488) && (pixel_index <= 3499)) || ((pixel_index >= 3503) && (pixel_index <= 3520)) || ((pixel_index >= 3523) && (pixel_index <= 3581)) || ((pixel_index >= 3584) && (pixel_index <= 3595)) || ((pixel_index >= 3599) && (pixel_index <= 3616)) || ((pixel_index >= 3619) && (pixel_index <= 3677)) || ((pixel_index >= 3680) && (pixel_index <= 3691)) || ((pixel_index >= 3694) && (pixel_index <= 3712)) || ((pixel_index >= 3715) && (pixel_index <= 3773)) || ((pixel_index >= 3776) && (pixel_index <= 3786)) || ((pixel_index >= 3790) && (pixel_index <= 3807)) || ((pixel_index >= 3811) && (pixel_index <= 3869)) || ((pixel_index >= 3872) && (pixel_index <= 3882)) || ((pixel_index >= 3886) && (pixel_index <= 3903)) || ((pixel_index >= 3907) && (pixel_index <= 3965)) || ((pixel_index >= 3968) && (pixel_index <= 3977)) || ((pixel_index >= 3981) && (pixel_index <= 3986)) || ((pixel_index >= 3988) && (pixel_index <= 3998)) || ((pixel_index >= 4002) && (pixel_index <= 4061)) || ((pixel_index >= 4064) && (pixel_index <= 4070)) || ((pixel_index >= 4077) && (pixel_index <= 4082)) || ((pixel_index >= 4086) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4157)) || ((pixel_index >= 4171) && (pixel_index <= 4178)) || ((pixel_index >= 4192) && (pixel_index <= 4253)) || ((pixel_index >= 4265) && (pixel_index <= 4276)) || (pixel_index >= 4286) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2156 || pixel_index == 3403 || pixel_index == 3598) oled_data = 16'b0101001010001010;
    else if (pixel_index == 3213 || pixel_index == 3502) oled_data = 16'b1010010100010100;
    else if (pixel_index == 3328) oled_data = 16'b1010011110010100;
    else oled_data = 0;
    end
    
    else if (freq>=1046 && freq<1108) //C6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1762)) || ((pixel_index >= 1772) && (pixel_index <= 1784)) || ((pixel_index >= 1795) && (pixel_index <= 1856)) || ((pixel_index >= 1870) && (pixel_index <= 1879)) || ((pixel_index >= 1891) && (pixel_index <= 1951)) || ((pixel_index >= 1956) && (pixel_index <= 1962)) || ((pixel_index >= 1967) && (pixel_index <= 1974)) || ((pixel_index >= 1978) && (pixel_index <= 1985)) || ((pixel_index >= 1987) && (pixel_index <= 2046)) || ((pixel_index >= 2051) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2069)) || ((pixel_index >= 2073) && (pixel_index <= 2141)) || ((pixel_index >= 2145) && (pixel_index <= 2157)) || ((pixel_index >= 2159) && (pixel_index <= 2164)) || ((pixel_index >= 2168) && (pixel_index <= 2237)) || ((pixel_index >= 2241) && (pixel_index <= 2260)) || ((pixel_index >= 2263) && (pixel_index <= 2332)) || ((pixel_index >= 2336) && (pixel_index <= 2355)) || ((pixel_index >= 2359) && (pixel_index <= 2428)) || ((pixel_index >= 2432) && (pixel_index <= 2451)) || ((pixel_index >= 2455) && (pixel_index <= 2524)) || ((pixel_index >= 2527) && (pixel_index <= 2547)) || ((pixel_index >= 2550) && (pixel_index <= 2619)) || ((pixel_index >= 2623) && (pixel_index <= 2642)) || ((pixel_index >= 2646) && (pixel_index <= 2715)) || ((pixel_index >= 2719) && (pixel_index <= 2738)) || ((pixel_index >= 2742) && (pixel_index <= 2811)) || ((pixel_index >= 2815) && (pixel_index <= 2834)) || pixel_index == 2838 || ((pixel_index >= 2849) && (pixel_index <= 2907)) || ((pixel_index >= 2911) && (pixel_index <= 2930)) || ((pixel_index >= 2946) && (pixel_index <= 3003)) || ((pixel_index >= 3007) && (pixel_index <= 3026)) || ((pixel_index >= 3032) && (pixel_index <= 3039)) || ((pixel_index >= 3043) && (pixel_index <= 3099)) || ((pixel_index >= 3103) && (pixel_index <= 3122)) || ((pixel_index >= 3126) && (pixel_index <= 3136)) || ((pixel_index >= 3140) && (pixel_index <= 3195)) || ((pixel_index >= 3199) && (pixel_index <= 3218)) || ((pixel_index >= 3222) && (pixel_index <= 3232)) || ((pixel_index >= 3236) && (pixel_index <= 3291)) || ((pixel_index >= 3295) && (pixel_index <= 3314)) || ((pixel_index >= 3318) && (pixel_index <= 3328)) || ((pixel_index >= 3332) && (pixel_index <= 3387)) || ((pixel_index >= 3391) && (pixel_index <= 3410)) || ((pixel_index >= 3414) && (pixel_index <= 3425)) || ((pixel_index >= 3428) && (pixel_index <= 3483)) || ((pixel_index >= 3487) && (pixel_index <= 3506)) || ((pixel_index >= 3510) && (pixel_index <= 3521)) || ((pixel_index >= 3524) && (pixel_index <= 3580)) || ((pixel_index >= 3584) && (pixel_index <= 3602)) || ((pixel_index >= 3606) && (pixel_index <= 3617)) || ((pixel_index >= 3620) && (pixel_index <= 3676)) || ((pixel_index >= 3680) && (pixel_index <= 3699)) || ((pixel_index >= 3702) && (pixel_index <= 3712)) || ((pixel_index >= 3716) && (pixel_index <= 3773)) || ((pixel_index >= 3777) && (pixel_index <= 3795)) || ((pixel_index >= 3799) && (pixel_index <= 3808)) || ((pixel_index >= 3812) && (pixel_index <= 3869)) || ((pixel_index >= 3874) && (pixel_index <= 3885)) || ((pixel_index >= 3887) && (pixel_index <= 3891)) || ((pixel_index >= 3895) && (pixel_index <= 3904)) || ((pixel_index >= 3908) && (pixel_index <= 3966)) || ((pixel_index >= 3971) && (pixel_index <= 3979)) || ((pixel_index >= 3983) && (pixel_index <= 3988)) || ((pixel_index >= 3992) && (pixel_index <= 3999)) || ((pixel_index >= 4003) && (pixel_index <= 4063)) || ((pixel_index >= 4069) && (pixel_index <= 4073)) || ((pixel_index >= 4079) && (pixel_index <= 4084)) || ((pixel_index >= 4089) && (pixel_index <= 4093)) || ((pixel_index >= 4098) && (pixel_index <= 4160)) || ((pixel_index >= 4174) && (pixel_index <= 4181)) || ((pixel_index >= 4193) && (pixel_index <= 4258)) || ((pixel_index >= 4267) && (pixel_index <= 4279)) || (pixel_index >= 4287) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2050 || pixel_index == 2839 || pixel_index == 3329 || pixel_index == 3907 || pixel_index == 4173) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2454) oled_data = 16'b0101010100001010;
    else oled_data = 0;
    end
    
    else if (freq>=1108 && freq<1174) //C#6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1389)) || ((pixel_index >= 1392) && (pixel_index <= 1395)) || ((pixel_index >= 1398) && (pixel_index <= 1485)) || ((pixel_index >= 1487) && (pixel_index <= 1491)) || ((pixel_index >= 1493) && (pixel_index <= 1581)) || ((pixel_index >= 1583) && (pixel_index <= 1587)) || ((pixel_index >= 1589) && (pixel_index <= 1676)) || ((pixel_index >= 1679) && (pixel_index <= 1682)) || ((pixel_index >= 1685) && (pixel_index <= 1755)) || ((pixel_index >= 1765) && (pixel_index <= 1772)) || ((pixel_index >= 1775) && (pixel_index <= 1778)) || ((pixel_index >= 1781) && (pixel_index <= 1791)) || ((pixel_index >= 1802) && (pixel_index <= 1849)) || ((pixel_index >= 1863) && (pixel_index <= 1866)) || ((pixel_index >= 1879) && (pixel_index <= 1886)) || ((pixel_index >= 1898) && (pixel_index <= 1944)) || ((pixel_index >= 1949) && (pixel_index <= 1955)) || ((pixel_index >= 1960) && (pixel_index <= 1964)) || ((pixel_index >= 1967) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 1981)) || ((pixel_index >= 1985) && (pixel_index <= 1992)) || ((pixel_index >= 1994) && (pixel_index <= 2039)) || ((pixel_index >= 2043) && (pixel_index <= 2053)) || ((pixel_index >= 2056) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2076)) || ((pixel_index >= 2080) && (pixel_index <= 2134)) || ((pixel_index >= 2138) && (pixel_index <= 2150)) || ((pixel_index >= 2152) && (pixel_index <= 2156)) || ((pixel_index >= 2159) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2171)) || ((pixel_index >= 2175) && (pixel_index <= 2230)) || ((pixel_index >= 2234) && (pixel_index <= 2252)) || ((pixel_index >= 2254) && (pixel_index <= 2258)) || ((pixel_index >= 2260) && (pixel_index <= 2267)) || ((pixel_index >= 2270) && (pixel_index <= 2325)) || ((pixel_index >= 2329) && (pixel_index <= 2348)) || ((pixel_index >= 2350) && (pixel_index <= 2354)) || ((pixel_index >= 2356) && (pixel_index <= 2362)) || ((pixel_index >= 2366) && (pixel_index <= 2421)) || ((pixel_index >= 2425) && (pixel_index <= 2441)) || ((pixel_index >= 2454) && (pixel_index <= 2458)) || ((pixel_index >= 2462) && (pixel_index <= 2516)) || ((pixel_index >= 2520) && (pixel_index <= 2537)) || ((pixel_index >= 2550) && (pixel_index <= 2554)) || ((pixel_index >= 2557) && (pixel_index <= 2612)) || ((pixel_index >= 2616) && (pixel_index <= 2635)) || ((pixel_index >= 2638) && (pixel_index <= 2641)) || ((pixel_index >= 2644) && (pixel_index <= 2650)) || ((pixel_index >= 2653) && (pixel_index <= 2708)) || ((pixel_index >= 2712) && (pixel_index <= 2731)) || ((pixel_index >= 2734) && (pixel_index <= 2737)) || ((pixel_index >= 2740) && (pixel_index <= 2745)) || ((pixel_index >= 2749) && (pixel_index <= 2804)) || ((pixel_index >= 2808) && (pixel_index <= 2827)) || ((pixel_index >= 2830) && (pixel_index <= 2833)) || ((pixel_index >= 2836) && (pixel_index <= 2841)) || ((pixel_index >= 2845) && (pixel_index <= 2846)) || ((pixel_index >= 2856) && (pixel_index <= 2900)) || ((pixel_index >= 2904) && (pixel_index <= 2923)) || ((pixel_index >= 2926) && (pixel_index <= 2929)) || ((pixel_index >= 2932) && (pixel_index <= 2937)) || ((pixel_index >= 2954) && (pixel_index <= 2996)) || ((pixel_index >= 3000) && (pixel_index <= 3019)) || ((pixel_index >= 3021) && (pixel_index <= 3025)) || ((pixel_index >= 3027) && (pixel_index <= 3033)) || ((pixel_index >= 3039) && (pixel_index <= 3046)) || ((pixel_index >= 3050) && (pixel_index <= 3092)) || ((pixel_index >= 3096) && (pixel_index <= 3129)) || ((pixel_index >= 3133) && (pixel_index <= 3143)) || ((pixel_index >= 3147) && (pixel_index <= 3188)) || ((pixel_index >= 3192) && (pixel_index <= 3225)) || ((pixel_index >= 3229) && (pixel_index <= 3239)) || ((pixel_index >= 3243) && (pixel_index <= 3284)) || ((pixel_index >= 3288) && (pixel_index <= 3321)) || ((pixel_index >= 3325) && (pixel_index <= 3336)) || ((pixel_index >= 3339) && (pixel_index <= 3380)) || ((pixel_index >= 3384) && (pixel_index <= 3417)) || ((pixel_index >= 3421) && (pixel_index <= 3432)) || ((pixel_index >= 3435) && (pixel_index <= 3476)) || ((pixel_index >= 3480) && (pixel_index <= 3513)) || ((pixel_index >= 3517) && (pixel_index <= 3528)) || ((pixel_index >= 3531) && (pixel_index <= 3573)) || ((pixel_index >= 3577) && (pixel_index <= 3610)) || ((pixel_index >= 3613) && (pixel_index <= 3624)) || ((pixel_index >= 3627) && (pixel_index <= 3669)) || ((pixel_index >= 3673) && (pixel_index <= 3706)) || ((pixel_index >= 3709) && (pixel_index <= 3720)) || ((pixel_index >= 3723) && (pixel_index <= 3765)) || ((pixel_index >= 3770) && (pixel_index <= 3802)) || ((pixel_index >= 3806) && (pixel_index <= 3815)) || ((pixel_index >= 3819) && (pixel_index <= 3862)) || ((pixel_index >= 3866) && (pixel_index <= 3878)) || ((pixel_index >= 3880) && (pixel_index <= 3898)) || ((pixel_index >= 3902) && (pixel_index <= 3911)) || ((pixel_index >= 3915) && (pixel_index <= 3959)) || ((pixel_index >= 3964) && (pixel_index <= 3972)) || ((pixel_index >= 3976) && (pixel_index <= 3995)) || ((pixel_index >= 3999) && (pixel_index <= 4006)) || ((pixel_index >= 4010) && (pixel_index <= 4056)) || ((pixel_index >= 4062) && (pixel_index <= 4066)) || ((pixel_index >= 4072) && (pixel_index <= 4091)) || ((pixel_index >= 4096) && (pixel_index <= 4100)) || ((pixel_index >= 4105) && (pixel_index <= 4153)) || ((pixel_index >= 4166) && (pixel_index <= 4188)) || ((pixel_index >= 4200) && (pixel_index <= 4251)) || ((pixel_index >= 4260) && (pixel_index <= 4286)) || (pixel_index >= 4294) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1397) oled_data = 16'b0000001010000000;
    else if (pixel_index == 1677 || pixel_index == 2164 || pixel_index == 2953) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2931) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=1174 && freq<1244) //D6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1755)) || ((pixel_index >= 1768) && (pixel_index <= 1786)) || ((pixel_index >= 1796) && (pixel_index <= 1851)) || ((pixel_index >= 1866) && (pixel_index <= 1880)) || ((pixel_index >= 1893) && (pixel_index <= 1947)) || ((pixel_index >= 1951) && (pixel_index <= 1957)) || ((pixel_index >= 1964) && (pixel_index <= 1975)) || ((pixel_index >= 1980) && (pixel_index <= 1987)) || ((pixel_index >= 1989) && (pixel_index <= 2043)) || ((pixel_index >= 2047) && (pixel_index <= 2056)) || ((pixel_index >= 2061) && (pixel_index <= 2070)) || ((pixel_index >= 2074) && (pixel_index <= 2139)) || ((pixel_index >= 2143) && (pixel_index <= 2153)) || ((pixel_index >= 2158) && (pixel_index <= 2166)) || ((pixel_index >= 2170) && (pixel_index <= 2235)) || ((pixel_index >= 2239) && (pixel_index <= 2250)) || ((pixel_index >= 2254) && (pixel_index <= 2261)) || ((pixel_index >= 2265) && (pixel_index <= 2331)) || ((pixel_index >= 2335) && (pixel_index <= 2347)) || ((pixel_index >= 2351) && (pixel_index <= 2357)) || ((pixel_index >= 2360) && (pixel_index <= 2427)) || ((pixel_index >= 2431) && (pixel_index <= 2443)) || ((pixel_index >= 2447) && (pixel_index <= 2452)) || ((pixel_index >= 2456) && (pixel_index <= 2523)) || ((pixel_index >= 2527) && (pixel_index <= 2540)) || ((pixel_index >= 2543) && (pixel_index <= 2548)) || ((pixel_index >= 2552) && (pixel_index <= 2619)) || ((pixel_index >= 2623) && (pixel_index <= 2636)) || ((pixel_index >= 2640) && (pixel_index <= 2644)) || ((pixel_index >= 2648) && (pixel_index <= 2715)) || ((pixel_index >= 2719) && (pixel_index <= 2732)) || ((pixel_index >= 2736) && (pixel_index <= 2740)) || ((pixel_index >= 2743) && (pixel_index <= 2811)) || ((pixel_index >= 2815) && (pixel_index <= 2828)) || ((pixel_index >= 2832) && (pixel_index <= 2836)) || ((pixel_index >= 2839) && (pixel_index <= 2840)) || ((pixel_index >= 2851) && (pixel_index <= 2907)) || ((pixel_index >= 2911) && (pixel_index <= 2924)) || ((pixel_index >= 2928) && (pixel_index <= 2932)) || ((pixel_index >= 2948) && (pixel_index <= 3003)) || ((pixel_index >= 3007) && (pixel_index <= 3020)) || ((pixel_index >= 3024) && (pixel_index <= 3028)) || ((pixel_index >= 3033) && (pixel_index <= 3040)) || ((pixel_index >= 3045) && (pixel_index <= 3099)) || ((pixel_index >= 3103) && (pixel_index <= 3116)) || ((pixel_index >= 3120) && (pixel_index <= 3124)) || ((pixel_index >= 3128) && (pixel_index <= 3137)) || ((pixel_index >= 3141) && (pixel_index <= 3195)) || ((pixel_index >= 3199) && (pixel_index <= 3212)) || ((pixel_index >= 3216) && (pixel_index <= 3220)) || ((pixel_index >= 3223) && (pixel_index <= 3234)) || ((pixel_index >= 3238) && (pixel_index <= 3291)) || ((pixel_index >= 3295) && (pixel_index <= 3308)) || ((pixel_index >= 3312) && (pixel_index <= 3316)) || ((pixel_index >= 3319) && (pixel_index <= 3330)) || ((pixel_index >= 3334) && (pixel_index <= 3387)) || ((pixel_index >= 3391) && (pixel_index <= 3404)) || ((pixel_index >= 3408) && (pixel_index <= 3412)) || ((pixel_index >= 3415) && (pixel_index <= 3426)) || ((pixel_index >= 3430) && (pixel_index <= 3483)) || ((pixel_index >= 3487) && (pixel_index <= 3499)) || ((pixel_index >= 3503) && (pixel_index <= 3508)) || ((pixel_index >= 3512) && (pixel_index <= 3522)) || ((pixel_index >= 3526) && (pixel_index <= 3579)) || ((pixel_index >= 3583) && (pixel_index <= 3595)) || ((pixel_index >= 3599) && (pixel_index <= 3604)) || ((pixel_index >= 3608) && (pixel_index <= 3618)) || ((pixel_index >= 3622) && (pixel_index <= 3675)) || ((pixel_index >= 3679) && (pixel_index <= 3691)) || ((pixel_index >= 3695) && (pixel_index <= 3700)) || ((pixel_index >= 3704) && (pixel_index <= 3714)) || ((pixel_index >= 3718) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3786)) || ((pixel_index >= 3790) && (pixel_index <= 3796)) || ((pixel_index >= 3800) && (pixel_index <= 3810)) || ((pixel_index >= 3813) && (pixel_index <= 3867)) || ((pixel_index >= 3871) && (pixel_index <= 3881)) || ((pixel_index >= 3885) && (pixel_index <= 3893)) || ((pixel_index >= 3897) && (pixel_index <= 3905)) || ((pixel_index >= 3909) && (pixel_index <= 3963)) || ((pixel_index >= 3967) && (pixel_index <= 3975)) || ((pixel_index >= 3980) && (pixel_index <= 3989)) || ((pixel_index >= 3993) && (pixel_index <= 4000)) || ((pixel_index >= 4004) && (pixel_index <= 4059)) || ((pixel_index >= 4063) && (pixel_index <= 4067)) || ((pixel_index >= 4075) && (pixel_index <= 4086)) || ((pixel_index >= 4091) && (pixel_index <= 4095)) || ((pixel_index >= 4100) && (pixel_index <= 4155)) || ((pixel_index >= 4170) && (pixel_index <= 4183)) || ((pixel_index >= 4195) && (pixel_index <= 4251)) || ((pixel_index >= 4263) && (pixel_index <= 4280)) || (pixel_index >= 4289) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 3127 || pixel_index == 3500 || pixel_index == 4068) oled_data = 16'b1010010100010100;
    else oled_data = 0;

    end
    
    else if (freq>=1244 && freq<1318) //Eb6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1290)) || ((pixel_index >= 1292) && (pixel_index <= 1386)) || ((pixel_index >= 1388) && (pixel_index <= 1482)) || ((pixel_index >= 1484) && (pixel_index <= 1578)) || ((pixel_index >= 1580) && (pixel_index <= 1674)) || ((pixel_index >= 1676) && (pixel_index <= 1750)) || ((pixel_index >= 1766) && (pixel_index <= 1770)) || ((pixel_index >= 1772) && (pixel_index <= 1791)) || ((pixel_index >= 1801) && (pixel_index <= 1846)) || ((pixel_index >= 1862) && (pixel_index <= 1866)) || ((pixel_index >= 1868) && (pixel_index <= 1869)) || ((pixel_index >= 1875) && (pixel_index <= 1885)) || ((pixel_index >= 1898) && (pixel_index <= 1942)) || ((pixel_index >= 1946) && (pixel_index <= 1962)) || pixel_index == 1964 || ((pixel_index >= 1967) && (pixel_index <= 1969)) || ((pixel_index >= 1972) && (pixel_index <= 1980)) || ((pixel_index >= 1985) && (pixel_index <= 1992)) || ((pixel_index >= 1994) && (pixel_index <= 2038)) || ((pixel_index >= 2042) && (pixel_index <= 2058)) || ((pixel_index >= 2061) && (pixel_index <= 2066)) || ((pixel_index >= 2069) && (pixel_index <= 2075)) || ((pixel_index >= 2079) && (pixel_index <= 2134)) || ((pixel_index >= 2138) && (pixel_index <= 2154)) || ((pixel_index >= 2156) && (pixel_index <= 2162)) || ((pixel_index >= 2165) && (pixel_index <= 2171)) || ((pixel_index >= 2174) && (pixel_index <= 2230)) || ((pixel_index >= 2234) && (pixel_index <= 2250)) || ((pixel_index >= 2252) && (pixel_index <= 2259)) || ((pixel_index >= 2261) && (pixel_index <= 2266)) || ((pixel_index >= 2270) && (pixel_index <= 2326)) || ((pixel_index >= 2330) && (pixel_index <= 2346)) || ((pixel_index >= 2348) && (pixel_index <= 2355)) || ((pixel_index >= 2358) && (pixel_index <= 2362)) || ((pixel_index >= 2365) && (pixel_index <= 2422)) || ((pixel_index >= 2426) && (pixel_index <= 2442)) || ((pixel_index >= 2444) && (pixel_index <= 2451)) || ((pixel_index >= 2454) && (pixel_index <= 2457)) || ((pixel_index >= 2461) && (pixel_index <= 2518)) || ((pixel_index >= 2522) && (pixel_index <= 2538)) || ((pixel_index >= 2540) && (pixel_index <= 2547)) || ((pixel_index >= 2549) && (pixel_index <= 2553)) || ((pixel_index >= 2557) && (pixel_index <= 2614)) || ((pixel_index >= 2618) && (pixel_index <= 2634)) || ((pixel_index >= 2636) && (pixel_index <= 2643)) || ((pixel_index >= 2645) && (pixel_index <= 2649)) || ((pixel_index >= 2652) && (pixel_index <= 2710)) || ((pixel_index >= 2714) && (pixel_index <= 2730)) || ((pixel_index >= 2732) && (pixel_index <= 2738)) || ((pixel_index >= 2741) && (pixel_index <= 2745)) || ((pixel_index >= 2748) && (pixel_index <= 2806)) || ((pixel_index >= 2810) && (pixel_index <= 2826)) || ((pixel_index >= 2829) && (pixel_index <= 2834)) || ((pixel_index >= 2837) && (pixel_index <= 2841)) || ((pixel_index >= 2844) && (pixel_index <= 2845)) || ((pixel_index >= 2856) && (pixel_index <= 2902)) || ((pixel_index >= 2916) && (pixel_index <= 2922)) || ((pixel_index >= 2927) && (pixel_index <= 2929)) || ((pixel_index >= 2932) && (pixel_index <= 2937)) || ((pixel_index >= 2953) && (pixel_index <= 2998)) || ((pixel_index >= 3012) && (pixel_index <= 3018)) || ((pixel_index >= 3020) && (pixel_index <= 3021)) || ((pixel_index >= 3027) && (pixel_index <= 3033)) || ((pixel_index >= 3038) && (pixel_index <= 3045)) || ((pixel_index >= 3050) && (pixel_index <= 3094)) || ((pixel_index >= 3098) && (pixel_index <= 3128)) || ((pixel_index >= 3132) && (pixel_index <= 3142)) || ((pixel_index >= 3146) && (pixel_index <= 3190)) || ((pixel_index >= 3194) && (pixel_index <= 3225)) || ((pixel_index >= 3228) && (pixel_index <= 3239)) || ((pixel_index >= 3242) && (pixel_index <= 3286)) || ((pixel_index >= 3290) && (pixel_index <= 3321)) || ((pixel_index >= 3324) && (pixel_index <= 3335)) || ((pixel_index >= 3339) && (pixel_index <= 3382)) || ((pixel_index >= 3386) && (pixel_index <= 3417)) || ((pixel_index >= 3420) && (pixel_index <= 3431)) || ((pixel_index >= 3435) && (pixel_index <= 3478)) || ((pixel_index >= 3482) && (pixel_index <= 3513)) || ((pixel_index >= 3516) && (pixel_index <= 3527)) || ((pixel_index >= 3531) && (pixel_index <= 3574)) || ((pixel_index >= 3578) && (pixel_index <= 3609)) || ((pixel_index >= 3613) && (pixel_index <= 3623)) || ((pixel_index >= 3627) && (pixel_index <= 3670)) || ((pixel_index >= 3674) && (pixel_index <= 3705)) || ((pixel_index >= 3709) && (pixel_index <= 3719)) || ((pixel_index >= 3723) && (pixel_index <= 3766)) || ((pixel_index >= 3770) && (pixel_index <= 3801)) || ((pixel_index >= 3805) && (pixel_index <= 3815)) || ((pixel_index >= 3818) && (pixel_index <= 3862)) || ((pixel_index >= 3866) && (pixel_index <= 3898)) || ((pixel_index >= 3902) && (pixel_index <= 3910)) || ((pixel_index >= 3914) && (pixel_index <= 3958)) || ((pixel_index >= 3962) && (pixel_index <= 3994)) || ((pixel_index >= 3998) && (pixel_index <= 4005)) || ((pixel_index >= 4009) && (pixel_index <= 4054)) || ((pixel_index >= 4058) && (pixel_index <= 4091)) || ((pixel_index >= 4096) && (pixel_index <= 4100)) || ((pixel_index >= 4105) && (pixel_index <= 4150)) || ((pixel_index >= 4166) && (pixel_index <= 4188)) || ((pixel_index >= 4200) && (pixel_index <= 4247)) || ((pixel_index >= 4262) && (pixel_index <= 4285)) || (pixel_index >= 4294) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1765 || pixel_index == 1861 || pixel_index == 1993 || pixel_index == 2855 || pixel_index == 3129) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2357 || pixel_index == 4199) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=1318 && freq<1396) //E6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1758)) || ((pixel_index >= 1773) && (pixel_index <= 1783)) || ((pixel_index >= 1794) && (pixel_index <= 1854)) || ((pixel_index >= 1869) && (pixel_index <= 1878)) || ((pixel_index >= 1890) && (pixel_index <= 1950)) || ((pixel_index >= 1953) && (pixel_index <= 1973)) || ((pixel_index >= 1977) && (pixel_index <= 1984)) || ((pixel_index >= 1986) && (pixel_index <= 2046)) || ((pixel_index >= 2049) && (pixel_index <= 2068)) || ((pixel_index >= 2072) && (pixel_index <= 2142)) || ((pixel_index >= 2145) && (pixel_index <= 2163)) || ((pixel_index >= 2167) && (pixel_index <= 2238)) || ((pixel_index >= 2241) && (pixel_index <= 2259)) || ((pixel_index >= 2262) && (pixel_index <= 2334)) || ((pixel_index >= 2337) && (pixel_index <= 2354)) || ((pixel_index >= 2358) && (pixel_index <= 2430)) || ((pixel_index >= 2433) && (pixel_index <= 2450)) || ((pixel_index >= 2454) && (pixel_index <= 2526)) || ((pixel_index >= 2529) && (pixel_index <= 2546)) || ((pixel_index >= 2549) && (pixel_index <= 2622)) || ((pixel_index >= 2625) && (pixel_index <= 2641)) || ((pixel_index >= 2645) && (pixel_index <= 2718)) || ((pixel_index >= 2721) && (pixel_index <= 2737)) || ((pixel_index >= 2741) && (pixel_index <= 2814)) || ((pixel_index >= 2817) && (pixel_index <= 2833)) || pixel_index == 2837 || ((pixel_index >= 2848) && (pixel_index <= 2910)) || ((pixel_index >= 2923) && (pixel_index <= 2929)) || ((pixel_index >= 2945) && (pixel_index <= 3006)) || ((pixel_index >= 3019) && (pixel_index <= 3025)) || ((pixel_index >= 3031) && (pixel_index <= 3038)) || ((pixel_index >= 3042) && (pixel_index <= 3102)) || ((pixel_index >= 3105) && (pixel_index <= 3121)) || ((pixel_index >= 3125) && (pixel_index <= 3135)) || ((pixel_index >= 3139) && (pixel_index <= 3198)) || ((pixel_index >= 3201) && (pixel_index <= 3217)) || ((pixel_index >= 3221) && (pixel_index <= 3231)) || ((pixel_index >= 3235) && (pixel_index <= 3294)) || ((pixel_index >= 3297) && (pixel_index <= 3313)) || ((pixel_index >= 3317) && (pixel_index <= 3328)) || ((pixel_index >= 3331) && (pixel_index <= 3390)) || ((pixel_index >= 3393) && (pixel_index <= 3409)) || ((pixel_index >= 3413) && (pixel_index <= 3424)) || ((pixel_index >= 3427) && (pixel_index <= 3486)) || ((pixel_index >= 3489) && (pixel_index <= 3505)) || ((pixel_index >= 3509) && (pixel_index <= 3520)) || ((pixel_index >= 3523) && (pixel_index <= 3582)) || ((pixel_index >= 3585) && (pixel_index <= 3601)) || ((pixel_index >= 3605) && (pixel_index <= 3616)) || ((pixel_index >= 3619) && (pixel_index <= 3678)) || ((pixel_index >= 3681) && (pixel_index <= 3698)) || ((pixel_index >= 3701) && (pixel_index <= 3711)) || ((pixel_index >= 3715) && (pixel_index <= 3774)) || ((pixel_index >= 3777) && (pixel_index <= 3794)) || ((pixel_index >= 3798) && (pixel_index <= 3807)) || ((pixel_index >= 3811) && (pixel_index <= 3870)) || ((pixel_index >= 3873) && (pixel_index <= 3890)) || ((pixel_index >= 3894) && (pixel_index <= 3903)) || ((pixel_index >= 3907) && (pixel_index <= 3966)) || ((pixel_index >= 3969) && (pixel_index <= 3987)) || ((pixel_index >= 3991) && (pixel_index <= 3998)) || ((pixel_index >= 4002) && (pixel_index <= 4062)) || ((pixel_index >= 4065) && (pixel_index <= 4083)) || ((pixel_index >= 4088) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4158)) || ((pixel_index >= 4173) && (pixel_index <= 4180)) || ((pixel_index >= 4192) && (pixel_index <= 4254)) || ((pixel_index >= 4269) && (pixel_index <= 4278)) || (pixel_index >= 4286) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2642 || pixel_index == 3906) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2838) oled_data = 16'b1010011110010100;
    else oled_data = 0;
    end
    
    else if (freq>=1396 && freq<1480) //F6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1758)) || ((pixel_index >= 1773) && (pixel_index <= 1783)) || ((pixel_index >= 1793) && (pixel_index <= 1854)) || ((pixel_index >= 1869) && (pixel_index <= 1877)) || ((pixel_index >= 1890) && (pixel_index <= 1950)) || ((pixel_index >= 1954) && (pixel_index <= 1972)) || ((pixel_index >= 1977) && (pixel_index <= 2046)) || ((pixel_index >= 2050) && (pixel_index <= 2067)) || ((pixel_index >= 2071) && (pixel_index <= 2142)) || ((pixel_index >= 2146) && (pixel_index <= 2163)) || ((pixel_index >= 2166) && (pixel_index <= 2238)) || ((pixel_index >= 2242) && (pixel_index <= 2258)) || ((pixel_index >= 2262) && (pixel_index <= 2334)) || ((pixel_index >= 2338) && (pixel_index <= 2354)) || ((pixel_index >= 2357) && (pixel_index <= 2430)) || ((pixel_index >= 2434) && (pixel_index <= 2449)) || ((pixel_index >= 2453) && (pixel_index <= 2526)) || ((pixel_index >= 2530) && (pixel_index <= 2545)) || ((pixel_index >= 2549) && (pixel_index <= 2622)) || ((pixel_index >= 2626) && (pixel_index <= 2641)) || ((pixel_index >= 2644) && (pixel_index <= 2718)) || ((pixel_index >= 2722) && (pixel_index <= 2737)) || ((pixel_index >= 2740) && (pixel_index <= 2814)) || ((pixel_index >= 2818) && (pixel_index <= 2833)) || ((pixel_index >= 2836) && (pixel_index <= 2837)) || ((pixel_index >= 2847) && (pixel_index <= 2910)) || ((pixel_index >= 2924) && (pixel_index <= 2928)) || ((pixel_index >= 2945) && (pixel_index <= 3006)) || ((pixel_index >= 3020) && (pixel_index <= 3024)) || ((pixel_index >= 3030) && (pixel_index <= 3037)) || ((pixel_index >= 3042) && (pixel_index <= 3102)) || ((pixel_index >= 3116) && (pixel_index <= 3120)) || ((pixel_index >= 3124) && (pixel_index <= 3134)) || ((pixel_index >= 3138) && (pixel_index <= 3198)) || ((pixel_index >= 3202) && (pixel_index <= 3216)) || ((pixel_index >= 3220) && (pixel_index <= 3231)) || ((pixel_index >= 3234) && (pixel_index <= 3294)) || ((pixel_index >= 3298) && (pixel_index <= 3313)) || ((pixel_index >= 3316) && (pixel_index <= 3327)) || ((pixel_index >= 3331) && (pixel_index <= 3390)) || ((pixel_index >= 3394) && (pixel_index <= 3409)) || ((pixel_index >= 3412) && (pixel_index <= 3423)) || ((pixel_index >= 3427) && (pixel_index <= 3486)) || ((pixel_index >= 3490) && (pixel_index <= 3505)) || ((pixel_index >= 3508) && (pixel_index <= 3519)) || ((pixel_index >= 3523) && (pixel_index <= 3582)) || ((pixel_index >= 3586) && (pixel_index <= 3601)) || ((pixel_index >= 3605) && (pixel_index <= 3615)) || ((pixel_index >= 3619) && (pixel_index <= 3678)) || ((pixel_index >= 3682) && (pixel_index <= 3697)) || ((pixel_index >= 3701) && (pixel_index <= 3711)) || ((pixel_index >= 3715) && (pixel_index <= 3774)) || ((pixel_index >= 3778) && (pixel_index <= 3793)) || ((pixel_index >= 3797) && (pixel_index <= 3806)) || ((pixel_index >= 3810) && (pixel_index <= 3870)) || ((pixel_index >= 3874) && (pixel_index <= 3890)) || ((pixel_index >= 3894) && (pixel_index <= 3902)) || ((pixel_index >= 3906) && (pixel_index <= 3966)) || ((pixel_index >= 3970) && (pixel_index <= 3986)) || ((pixel_index >= 3990) && (pixel_index <= 3997)) || ((pixel_index >= 4001) && (pixel_index <= 4062)) || ((pixel_index >= 4066) && (pixel_index <= 4083)) || ((pixel_index >= 4088) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4158)) || ((pixel_index >= 4162) && (pixel_index <= 4180)) || ((pixel_index >= 4191) && (pixel_index <= 4254)) || ((pixel_index >= 4258) && (pixel_index <= 4277)) || (pixel_index >= 4286) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2929) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=1480 && freq<1568) //F#6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1387)) || ((pixel_index >= 1390) && (pixel_index <= 1393)) || ((pixel_index >= 1396) && (pixel_index <= 1483)) || ((pixel_index >= 1486) && (pixel_index <= 1489)) || ((pixel_index >= 1492) && (pixel_index <= 1579)) || ((pixel_index >= 1582) && (pixel_index <= 1585)) || ((pixel_index >= 1588) && (pixel_index <= 1675)) || ((pixel_index >= 1678) && (pixel_index <= 1681)) || ((pixel_index >= 1684) && (pixel_index <= 1751)) || ((pixel_index >= 1766) && (pixel_index <= 1771)) || ((pixel_index >= 1773) && (pixel_index <= 1777)) || ((pixel_index >= 1779) && (pixel_index <= 1790)) || ((pixel_index >= 1800) && (pixel_index <= 1847)) || ((pixel_index >= 1862) && (pixel_index <= 1864)) || ((pixel_index >= 1878) && (pixel_index <= 1884)) || ((pixel_index >= 1897) && (pixel_index <= 1943)) || ((pixel_index >= 1947) && (pixel_index <= 1962)) || ((pixel_index >= 1965) && (pixel_index <= 1968)) || ((pixel_index >= 1971) && (pixel_index <= 1979)) || ((pixel_index >= 1984) && (pixel_index <= 1991)) || ((pixel_index >= 1993) && (pixel_index <= 2039)) || ((pixel_index >= 2043) && (pixel_index <= 2058)) || ((pixel_index >= 2061) && (pixel_index <= 2064)) || ((pixel_index >= 2067) && (pixel_index <= 2074)) || ((pixel_index >= 2078) && (pixel_index <= 2135)) || ((pixel_index >= 2139) && (pixel_index <= 2154)) || ((pixel_index >= 2157) && (pixel_index <= 2160)) || ((pixel_index >= 2163) && (pixel_index <= 2170)) || ((pixel_index >= 2174) && (pixel_index <= 2231)) || ((pixel_index >= 2235) && (pixel_index <= 2250)) || ((pixel_index >= 2253) && (pixel_index <= 2256)) || ((pixel_index >= 2259) && (pixel_index <= 2265)) || ((pixel_index >= 2269) && (pixel_index <= 2327)) || ((pixel_index >= 2331) && (pixel_index <= 2346)) || ((pixel_index >= 2349) && (pixel_index <= 2352)) || ((pixel_index >= 2355) && (pixel_index <= 2361)) || ((pixel_index >= 2364) && (pixel_index <= 2423)) || ((pixel_index >= 2427) && (pixel_index <= 2440)) || ((pixel_index >= 2453) && (pixel_index <= 2456)) || ((pixel_index >= 2460) && (pixel_index <= 2519)) || ((pixel_index >= 2523) && (pixel_index <= 2535)) || ((pixel_index >= 2549) && (pixel_index <= 2552)) || ((pixel_index >= 2556) && (pixel_index <= 2615)) || ((pixel_index >= 2619) && (pixel_index <= 2634)) || ((pixel_index >= 2636) && (pixel_index <= 2640)) || ((pixel_index >= 2642) && (pixel_index <= 2648)) || ((pixel_index >= 2652) && (pixel_index <= 2711)) || ((pixel_index >= 2715) && (pixel_index <= 2729)) || ((pixel_index >= 2732) && (pixel_index <= 2735)) || ((pixel_index >= 2738) && (pixel_index <= 2744)) || ((pixel_index >= 2747) && (pixel_index <= 2807)) || ((pixel_index >= 2811) && (pixel_index <= 2825)) || ((pixel_index >= 2828) && (pixel_index <= 2831)) || ((pixel_index >= 2834) && (pixel_index <= 2840)) || ((pixel_index >= 2843) && (pixel_index <= 2844)) || ((pixel_index >= 2855) && (pixel_index <= 2903)) || ((pixel_index >= 2917) && (pixel_index <= 2921)) || ((pixel_index >= 2924) && (pixel_index <= 2927)) || ((pixel_index >= 2930) && (pixel_index <= 2936)) || ((pixel_index >= 2952) && (pixel_index <= 2999)) || ((pixel_index >= 3013) && (pixel_index <= 3017)) || ((pixel_index >= 3020) && (pixel_index <= 3023)) || ((pixel_index >= 3026) && (pixel_index <= 3032)) || ((pixel_index >= 3037) && (pixel_index <= 3044)) || ((pixel_index >= 3049) && (pixel_index <= 3095)) || ((pixel_index >= 3109) && (pixel_index <= 3128)) || ((pixel_index >= 3131) && (pixel_index <= 3141)) || ((pixel_index >= 3145) && (pixel_index <= 3191)) || ((pixel_index >= 3195) && (pixel_index <= 3224)) || ((pixel_index >= 3227) && (pixel_index <= 3238)) || ((pixel_index >= 3242) && (pixel_index <= 3287)) || ((pixel_index >= 3291) && (pixel_index <= 3320)) || ((pixel_index >= 3323) && (pixel_index <= 3334)) || ((pixel_index >= 3338) && (pixel_index <= 3383)) || ((pixel_index >= 3387) && (pixel_index <= 3416)) || ((pixel_index >= 3419) && (pixel_index <= 3430)) || ((pixel_index >= 3434) && (pixel_index <= 3479)) || ((pixel_index >= 3483) && (pixel_index <= 3512)) || ((pixel_index >= 3515) && (pixel_index <= 3526)) || ((pixel_index >= 3530) && (pixel_index <= 3575)) || ((pixel_index >= 3579) && (pixel_index <= 3608)) || ((pixel_index >= 3612) && (pixel_index <= 3622)) || ((pixel_index >= 3626) && (pixel_index <= 3671)) || ((pixel_index >= 3675) && (pixel_index <= 3704)) || ((pixel_index >= 3708) && (pixel_index <= 3718)) || ((pixel_index >= 3722) && (pixel_index <= 3767)) || ((pixel_index >= 3771) && (pixel_index <= 3800)) || ((pixel_index >= 3804) && (pixel_index <= 3814)) || ((pixel_index >= 3817) && (pixel_index <= 3863)) || ((pixel_index >= 3867) && (pixel_index <= 3897)) || ((pixel_index >= 3901) && (pixel_index <= 3909)) || ((pixel_index >= 3913) && (pixel_index <= 3959)) || ((pixel_index >= 3963) && (pixel_index <= 3993)) || ((pixel_index >= 3997) && (pixel_index <= 4004)) || ((pixel_index >= 4008) && (pixel_index <= 4055)) || ((pixel_index >= 4059) && (pixel_index <= 4090)) || ((pixel_index >= 4095) && (pixel_index <= 4099)) || ((pixel_index >= 4104) && (pixel_index <= 4151)) || ((pixel_index >= 4155) && (pixel_index <= 4187)) || ((pixel_index >= 4199) && (pixel_index <= 4247)) || ((pixel_index >= 4251) && (pixel_index <= 4284)) || (pixel_index >= 4293) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1963 || pixel_index == 2854) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2173 || pixel_index == 2651) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2536) oled_data = 16'b1010011110010100;
    else oled_data = 0;
    end
    
    else if (freq>=1568 && freq<1661) //G6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1761)) || ((pixel_index >= 1772) && (pixel_index <= 1786)) || ((pixel_index >= 1797) && (pixel_index <= 1855)) || ((pixel_index >= 1870) && (pixel_index <= 1881)) || ((pixel_index >= 1893) && (pixel_index <= 1949)) || ((pixel_index >= 1955) && (pixel_index <= 1962)) || ((pixel_index >= 1967) && (pixel_index <= 1976)) || ((pixel_index >= 1980) && (pixel_index <= 1987)) || ((pixel_index >= 1989) && (pixel_index <= 2044)) || ((pixel_index >= 2049) && (pixel_index <= 2060)) || ((pixel_index >= 2063) && (pixel_index <= 2071)) || ((pixel_index >= 2075) && (pixel_index <= 2140)) || ((pixel_index >= 2144) && (pixel_index <= 2166)) || ((pixel_index >= 2170) && (pixel_index <= 2235)) || ((pixel_index >= 2239) && (pixel_index <= 2262)) || ((pixel_index >= 2265) && (pixel_index <= 2330)) || ((pixel_index >= 2334) && (pixel_index <= 2357)) || ((pixel_index >= 2361) && (pixel_index <= 2426)) || ((pixel_index >= 2430) && (pixel_index <= 2453)) || ((pixel_index >= 2457) && (pixel_index <= 2522)) || ((pixel_index >= 2525) && (pixel_index <= 2549)) || ((pixel_index >= 2552) && (pixel_index <= 2617)) || ((pixel_index >= 2621) && (pixel_index <= 2644)) || ((pixel_index >= 2648) && (pixel_index <= 2713)) || ((pixel_index >= 2717) && (pixel_index <= 2740)) || ((pixel_index >= 2744) && (pixel_index <= 2809)) || ((pixel_index >= 2813) && (pixel_index <= 2836)) || pixel_index == 2840 || ((pixel_index >= 2851) && (pixel_index <= 2905)) || ((pixel_index >= 2909) && (pixel_index <= 2916)) || ((pixel_index >= 2927) && (pixel_index <= 2932)) || ((pixel_index >= 2948) && (pixel_index <= 3001)) || ((pixel_index >= 3005) && (pixel_index <= 3012)) || ((pixel_index >= 3023) && (pixel_index <= 3028)) || ((pixel_index >= 3034) && (pixel_index <= 3041)) || ((pixel_index >= 3045) && (pixel_index <= 3097)) || ((pixel_index >= 3101) && (pixel_index <= 3108)) || ((pixel_index >= 3119) && (pixel_index <= 3124)) || ((pixel_index >= 3128) && (pixel_index <= 3138)) || ((pixel_index >= 3142) && (pixel_index <= 3193)) || ((pixel_index >= 3197) && (pixel_index <= 3212)) || ((pixel_index >= 3215) && (pixel_index <= 3220)) || ((pixel_index >= 3224) && (pixel_index <= 3234)) || ((pixel_index >= 3238) && (pixel_index <= 3289)) || ((pixel_index >= 3293) && (pixel_index <= 3308)) || ((pixel_index >= 3311) && (pixel_index <= 3316)) || ((pixel_index >= 3320) && (pixel_index <= 3330)) || ((pixel_index >= 3334) && (pixel_index <= 3385)) || ((pixel_index >= 3389) && (pixel_index <= 3404)) || ((pixel_index >= 3407) && (pixel_index <= 3412)) || ((pixel_index >= 3416) && (pixel_index <= 3427)) || ((pixel_index >= 3430) && (pixel_index <= 3482)) || ((pixel_index >= 3486) && (pixel_index <= 3500)) || ((pixel_index >= 3503) && (pixel_index <= 3508)) || ((pixel_index >= 3512) && (pixel_index <= 3523)) || ((pixel_index >= 3526) && (pixel_index <= 3578)) || ((pixel_index >= 3582) && (pixel_index <= 3596)) || ((pixel_index >= 3599) && (pixel_index <= 3604)) || ((pixel_index >= 3608) && (pixel_index <= 3619)) || ((pixel_index >= 3622) && (pixel_index <= 3674)) || ((pixel_index >= 3679) && (pixel_index <= 3692)) || ((pixel_index >= 3695) && (pixel_index <= 3701)) || ((pixel_index >= 3704) && (pixel_index <= 3714)) || ((pixel_index >= 3718) && (pixel_index <= 3771)) || ((pixel_index >= 3775) && (pixel_index <= 3788)) || ((pixel_index >= 3791) && (pixel_index <= 3797)) || ((pixel_index >= 3801) && (pixel_index <= 3810)) || ((pixel_index >= 3814) && (pixel_index <= 3868)) || ((pixel_index >= 3872) && (pixel_index <= 3884)) || ((pixel_index >= 3887) && (pixel_index <= 3893)) || ((pixel_index >= 3897) && (pixel_index <= 3906)) || ((pixel_index >= 3909) && (pixel_index <= 3964)) || ((pixel_index >= 3970) && (pixel_index <= 3979)) || ((pixel_index >= 3983) && (pixel_index <= 3990)) || ((pixel_index >= 3994) && (pixel_index <= 4001)) || ((pixel_index >= 4005) && (pixel_index <= 4061)) || ((pixel_index >= 4068) && (pixel_index <= 4073)) || ((pixel_index >= 4079) && (pixel_index <= 4086)) || ((pixel_index >= 4091) && (pixel_index <= 4095)) || ((pixel_index >= 4100) && (pixel_index <= 4159)) || ((pixel_index >= 4174) && (pixel_index <= 4183)) || ((pixel_index >= 4195) && (pixel_index <= 4257)) || ((pixel_index >= 4267) && (pixel_index <= 4281)) || (pixel_index >= 4289) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2456 || pixel_index == 2841) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2926 || pixel_index == 3331 || pixel_index == 3485 || pixel_index == 3678) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=1661 && freq<1760) //Ab6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1291)) || ((pixel_index >= 1294) && (pixel_index <= 1387)) || ((pixel_index >= 1390) && (pixel_index <= 1483)) || ((pixel_index >= 1486) && (pixel_index <= 1579)) || ((pixel_index >= 1582) && (pixel_index <= 1675)) || ((pixel_index >= 1678) && (pixel_index <= 1755)) || ((pixel_index >= 1759) && (pixel_index <= 1771)) || ((pixel_index >= 1774) && (pixel_index <= 1792)) || ((pixel_index >= 1803) && (pixel_index <= 1851)) || ((pixel_index >= 1856) && (pixel_index <= 1867)) || pixel_index == 1870 || ((pixel_index >= 1877) && (pixel_index <= 1887)) || ((pixel_index >= 1899) && (pixel_index <= 1946)) || ((pixel_index >= 1952) && (pixel_index <= 1963)) || ((pixel_index >= 1968) && (pixel_index <= 1970)) || ((pixel_index >= 1974) && (pixel_index <= 1982)) || ((pixel_index >= 1986) && (pixel_index <= 1993)) || ((pixel_index >= 1995) && (pixel_index <= 2042)) || pixel_index == 2045 || ((pixel_index >= 2049) && (pixel_index <= 2059)) || ((pixel_index >= 2063) && (pixel_index <= 2067)) || ((pixel_index >= 2070) && (pixel_index <= 2077)) || ((pixel_index >= 2081) && (pixel_index <= 2138)) || pixel_index == 2141 || ((pixel_index >= 2145) && (pixel_index <= 2155)) || ((pixel_index >= 2158) && (pixel_index <= 2164)) || ((pixel_index >= 2167) && (pixel_index <= 2172)) || ((pixel_index >= 2176) && (pixel_index <= 2233)) || ((pixel_index >= 2237) && (pixel_index <= 2238)) || ((pixel_index >= 2241) && (pixel_index <= 2251)) || ((pixel_index >= 2254) && (pixel_index <= 2260)) || ((pixel_index >= 2263) && (pixel_index <= 2268)) || ((pixel_index >= 2271) && (pixel_index <= 2329)) || ((pixel_index >= 2332) && (pixel_index <= 2334)) || ((pixel_index >= 2338) && (pixel_index <= 2347)) || ((pixel_index >= 2350) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2363)) || ((pixel_index >= 2367) && (pixel_index <= 2424)) || ((pixel_index >= 2428) && (pixel_index <= 2430)) || ((pixel_index >= 2434) && (pixel_index <= 2443)) || ((pixel_index >= 2446) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2459)) || ((pixel_index >= 2463) && (pixel_index <= 2520)) || ((pixel_index >= 2524) && (pixel_index <= 2527)) || ((pixel_index >= 2530) && (pixel_index <= 2539)) || ((pixel_index >= 2542) && (pixel_index <= 2548)) || ((pixel_index >= 2551) && (pixel_index <= 2555)) || ((pixel_index >= 2558) && (pixel_index <= 2616)) || ((pixel_index >= 2619) && (pixel_index <= 2623)) || ((pixel_index >= 2627) && (pixel_index <= 2635)) || ((pixel_index >= 2638) && (pixel_index <= 2644)) || ((pixel_index >= 2647) && (pixel_index <= 2650)) || ((pixel_index >= 2654) && (pixel_index <= 2711)) || ((pixel_index >= 2715) && (pixel_index <= 2719)) || ((pixel_index >= 2723) && (pixel_index <= 2731)) || ((pixel_index >= 2734) && (pixel_index <= 2740)) || ((pixel_index >= 2743) && (pixel_index <= 2746)) || ((pixel_index >= 2750) && (pixel_index <= 2807)) || ((pixel_index >= 2810) && (pixel_index <= 2816)) || ((pixel_index >= 2820) && (pixel_index <= 2827)) || ((pixel_index >= 2831) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2842)) || pixel_index == 2846 || ((pixel_index >= 2857) && (pixel_index <= 2903)) || ((pixel_index >= 2906) && (pixel_index <= 2912)) || ((pixel_index >= 2916) && (pixel_index <= 2923)) || ((pixel_index >= 2928) && (pixel_index <= 2930)) || ((pixel_index >= 2934) && (pixel_index <= 2938)) || ((pixel_index >= 2954) && (pixel_index <= 2998)) || ((pixel_index >= 3002) && (pixel_index <= 3009)) || ((pixel_index >= 3012) && (pixel_index <= 3019)) || pixel_index == 3022 || ((pixel_index >= 3029) && (pixel_index <= 3034)) || ((pixel_index >= 3040) && (pixel_index <= 3047)) || ((pixel_index >= 3051) && (pixel_index <= 3094)) || ((pixel_index >= 3097) && (pixel_index <= 3105)) || ((pixel_index >= 3109) && (pixel_index <= 3130)) || ((pixel_index >= 3134) && (pixel_index <= 3144)) || ((pixel_index >= 3148) && (pixel_index <= 3190)) || ((pixel_index >= 3193) && (pixel_index <= 3201)) || ((pixel_index >= 3205) && (pixel_index <= 3226)) || ((pixel_index >= 3230) && (pixel_index <= 3240)) || ((pixel_index >= 3244) && (pixel_index <= 3285)) || ((pixel_index >= 3289) && (pixel_index <= 3298)) || ((pixel_index >= 3301) && (pixel_index <= 3322)) || ((pixel_index >= 3326) && (pixel_index <= 3337)) || ((pixel_index >= 3340) && (pixel_index <= 3381)) || ((pixel_index >= 3398) && (pixel_index <= 3418)) || ((pixel_index >= 3422) && (pixel_index <= 3433)) || ((pixel_index >= 3436) && (pixel_index <= 3476)) || ((pixel_index >= 3494) && (pixel_index <= 3514)) || ((pixel_index >= 3518) && (pixel_index <= 3529)) || ((pixel_index >= 3532) && (pixel_index <= 3572)) || ((pixel_index >= 3576) && (pixel_index <= 3587)) || ((pixel_index >= 3590) && (pixel_index <= 3610)) || ((pixel_index >= 3614) && (pixel_index <= 3625)) || ((pixel_index >= 3628) && (pixel_index <= 3668)) || ((pixel_index >= 3671) && (pixel_index <= 3683)) || ((pixel_index >= 3687) && (pixel_index <= 3707)) || ((pixel_index >= 3710) && (pixel_index <= 3720)) || ((pixel_index >= 3724) && (pixel_index <= 3763)) || ((pixel_index >= 3767) && (pixel_index <= 3779)) || ((pixel_index >= 3783) && (pixel_index <= 3803)) || ((pixel_index >= 3807) && (pixel_index <= 3816)) || ((pixel_index >= 3820) && (pixel_index <= 3859)) || ((pixel_index >= 3863) && (pixel_index <= 3876)) || ((pixel_index >= 3880) && (pixel_index <= 3899)) || ((pixel_index >= 3903) && (pixel_index <= 3912)) || ((pixel_index >= 3916) && (pixel_index <= 3955)) || ((pixel_index >= 3958) && (pixel_index <= 3972)) || ((pixel_index >= 3976) && (pixel_index <= 3996)) || ((pixel_index >= 4000) && (pixel_index <= 4007)) || ((pixel_index >= 4011) && (pixel_index <= 4050)) || ((pixel_index >= 4054) && (pixel_index <= 4068)) || ((pixel_index >= 4072) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4101)) || ((pixel_index >= 4106) && (pixel_index <= 4146)) || ((pixel_index >= 4150) && (pixel_index <= 4165)) || ((pixel_index >= 4169) && (pixel_index <= 4189)) || ((pixel_index >= 4201) && (pixel_index <= 4242)) || ((pixel_index >= 4245) && (pixel_index <= 4261)) || ((pixel_index >= 4265) && (pixel_index <= 4287)) || (pixel_index >= 4295) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1971 || pixel_index == 2847) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2651 || pixel_index == 3915 || pixel_index == 4069) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2819) oled_data = 16'b0101010100001010;
    else oled_data = 0;
    end
    
    else if (freq>=1760 && freq<1864) //A6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1762)) || ((pixel_index >= 1767) && (pixel_index <= 1785)) || ((pixel_index >= 1795) && (pixel_index <= 1858)) || ((pixel_index >= 1863) && (pixel_index <= 1879)) || ((pixel_index >= 1892) && (pixel_index <= 1954)) || ((pixel_index >= 1960) && (pixel_index <= 1974)) || ((pixel_index >= 1979) && (pixel_index <= 1986)) || ((pixel_index >= 1988) && (pixel_index <= 2049)) || ((pixel_index >= 2056) && (pixel_index <= 2069)) || ((pixel_index >= 2074) && (pixel_index <= 2145)) || ((pixel_index >= 2148) && (pixel_index <= 2149)) || ((pixel_index >= 2152) && (pixel_index <= 2165)) || ((pixel_index >= 2169) && (pixel_index <= 2241)) || ((pixel_index >= 2244) && (pixel_index <= 2245)) || ((pixel_index >= 2249) && (pixel_index <= 2260)) || ((pixel_index >= 2264) && (pixel_index <= 2336)) || ((pixel_index >= 2340) && (pixel_index <= 2341)) || ((pixel_index >= 2345) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2432)) || ((pixel_index >= 2435) && (pixel_index <= 2438)) || ((pixel_index >= 2441) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2527)) || ((pixel_index >= 2531) && (pixel_index <= 2534)) || ((pixel_index >= 2538) && (pixel_index <= 2547)) || ((pixel_index >= 2551) && (pixel_index <= 2623)) || ((pixel_index >= 2627) && (pixel_index <= 2630)) || ((pixel_index >= 2634) && (pixel_index <= 2643)) || ((pixel_index >= 2647) && (pixel_index <= 2719)) || ((pixel_index >= 2722) && (pixel_index <= 2727)) || ((pixel_index >= 2731) && (pixel_index <= 2739)) || ((pixel_index >= 2742) && (pixel_index <= 2814)) || ((pixel_index >= 2818) && (pixel_index <= 2823)) || ((pixel_index >= 2827) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2839)) || ((pixel_index >= 2850) && (pixel_index <= 2910)) || ((pixel_index >= 2914) && (pixel_index <= 2920)) || ((pixel_index >= 2923) && (pixel_index <= 2931)) || ((pixel_index >= 2947) && (pixel_index <= 3006)) || ((pixel_index >= 3009) && (pixel_index <= 3016)) || ((pixel_index >= 3020) && (pixel_index <= 3027)) || ((pixel_index >= 3033) && (pixel_index <= 3039)) || ((pixel_index >= 3044) && (pixel_index <= 3101)) || ((pixel_index >= 3105) && (pixel_index <= 3112)) || ((pixel_index >= 3116) && (pixel_index <= 3123)) || ((pixel_index >= 3127) && (pixel_index <= 3136)) || ((pixel_index >= 3140) && (pixel_index <= 3197)) || ((pixel_index >= 3201) && (pixel_index <= 3209)) || ((pixel_index >= 3212) && (pixel_index <= 3219)) || ((pixel_index >= 3222) && (pixel_index <= 3233)) || ((pixel_index >= 3237) && (pixel_index <= 3293)) || ((pixel_index >= 3296) && (pixel_index <= 3305)) || ((pixel_index >= 3309) && (pixel_index <= 3315)) || ((pixel_index >= 3318) && (pixel_index <= 3329)) || ((pixel_index >= 3333) && (pixel_index <= 3388)) || ((pixel_index >= 3405) && (pixel_index <= 3411)) || ((pixel_index >= 3414) && (pixel_index <= 3425)) || ((pixel_index >= 3429) && (pixel_index <= 3484)) || ((pixel_index >= 3501) && (pixel_index <= 3507)) || ((pixel_index >= 3511) && (pixel_index <= 3521)) || ((pixel_index >= 3525) && (pixel_index <= 3579)) || ((pixel_index >= 3583) && (pixel_index <= 3594)) || ((pixel_index >= 3598) && (pixel_index <= 3603)) || ((pixel_index >= 3607) && (pixel_index <= 3617)) || ((pixel_index >= 3621) && (pixel_index <= 3675)) || ((pixel_index >= 3679) && (pixel_index <= 3690)) || ((pixel_index >= 3694) && (pixel_index <= 3699)) || ((pixel_index >= 3703) && (pixel_index <= 3713)) || ((pixel_index >= 3717) && (pixel_index <= 3771)) || ((pixel_index >= 3774) && (pixel_index <= 3787)) || ((pixel_index >= 3791) && (pixel_index <= 3796)) || ((pixel_index >= 3799) && (pixel_index <= 3809)) || ((pixel_index >= 3813) && (pixel_index <= 3866)) || ((pixel_index >= 3870) && (pixel_index <= 3883)) || ((pixel_index >= 3887) && (pixel_index <= 3892)) || ((pixel_index >= 3896) && (pixel_index <= 3904)) || ((pixel_index >= 3908) && (pixel_index <= 3962)) || ((pixel_index >= 3966) && (pixel_index <= 3980)) || ((pixel_index >= 3983) && (pixel_index <= 3988)) || ((pixel_index >= 3992) && (pixel_index <= 3999)) || ((pixel_index >= 4004) && (pixel_index <= 4058)) || ((pixel_index >= 4061) && (pixel_index <= 4076)) || ((pixel_index >= 4080) && (pixel_index <= 4085)) || ((pixel_index >= 4090) && (pixel_index <= 4094)) || ((pixel_index >= 4099) && (pixel_index <= 4153)) || ((pixel_index >= 4157) && (pixel_index <= 4172)) || ((pixel_index >= 4176) && (pixel_index <= 4182)) || ((pixel_index >= 4194) && (pixel_index <= 4249)) || ((pixel_index >= 4253) && (pixel_index <= 4269)) || ((pixel_index >= 4272) && (pixel_index <= 4279)) || (pixel_index >= 4288) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2528 || pixel_index == 2631 || pixel_index == 3032 || pixel_index == 3200 || pixel_index == 3812) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
    
    else if (freq>=1864 && freq<1975) //Bb6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1290)) || ((pixel_index >= 1293) && (pixel_index <= 1386)) || ((pixel_index >= 1389) && (pixel_index <= 1482)) || ((pixel_index >= 1485) && (pixel_index <= 1578)) || ((pixel_index >= 1581) && (pixel_index <= 1674)) || ((pixel_index >= 1677) && (pixel_index <= 1749)) || ((pixel_index >= 1762) && (pixel_index <= 1770)) || ((pixel_index >= 1773) && (pixel_index <= 1792)) || ((pixel_index >= 1802) && (pixel_index <= 1845)) || ((pixel_index >= 1859) && (pixel_index <= 1866)) || ((pixel_index >= 1869) && (pixel_index <= 1870)) || ((pixel_index >= 1876) && (pixel_index <= 1886)) || ((pixel_index >= 1899) && (pixel_index <= 1941)) || ((pixel_index >= 1945) && (pixel_index <= 1951)) || ((pixel_index >= 1956) && (pixel_index <= 1962)) || ((pixel_index >= 1968) && (pixel_index <= 1970)) || ((pixel_index >= 1973) && (pixel_index <= 1981)) || ((pixel_index >= 1986) && (pixel_index <= 2037)) || ((pixel_index >= 2041) && (pixel_index <= 2048)) || ((pixel_index >= 2053) && (pixel_index <= 2058)) || ((pixel_index >= 2062) && (pixel_index <= 2067)) || ((pixel_index >= 2070) && (pixel_index <= 2076)) || ((pixel_index >= 2080) && (pixel_index <= 2133)) || ((pixel_index >= 2137) && (pixel_index <= 2145)) || ((pixel_index >= 2149) && (pixel_index <= 2154)) || ((pixel_index >= 2157) && (pixel_index <= 2163)) || ((pixel_index >= 2166) && (pixel_index <= 2172)) || ((pixel_index >= 2175) && (pixel_index <= 2229)) || ((pixel_index >= 2233) && (pixel_index <= 2241)) || ((pixel_index >= 2245) && (pixel_index <= 2250)) || ((pixel_index >= 2253) && (pixel_index <= 2260)) || ((pixel_index >= 2262) && (pixel_index <= 2267)) || ((pixel_index >= 2271) && (pixel_index <= 2325)) || ((pixel_index >= 2329) && (pixel_index <= 2338)) || ((pixel_index >= 2341) && (pixel_index <= 2346)) || ((pixel_index >= 2349) && (pixel_index <= 2356)) || ((pixel_index >= 2359) && (pixel_index <= 2363)) || ((pixel_index >= 2366) && (pixel_index <= 2421)) || ((pixel_index >= 2425) && (pixel_index <= 2434)) || ((pixel_index >= 2437) && (pixel_index <= 2442)) || ((pixel_index >= 2445) && (pixel_index <= 2452)) || ((pixel_index >= 2455) && (pixel_index <= 2458)) || ((pixel_index >= 2462) && (pixel_index <= 2517)) || ((pixel_index >= 2521) && (pixel_index <= 2529)) || ((pixel_index >= 2533) && (pixel_index <= 2538)) || ((pixel_index >= 2541) && (pixel_index <= 2548)) || ((pixel_index >= 2550) && (pixel_index <= 2554)) || ((pixel_index >= 2558) && (pixel_index <= 2613)) || ((pixel_index >= 2617) && (pixel_index <= 2625)) || ((pixel_index >= 2629) && (pixel_index <= 2634)) || ((pixel_index >= 2637) && (pixel_index <= 2644)) || ((pixel_index >= 2646) && (pixel_index <= 2650)) || ((pixel_index >= 2653) && (pixel_index <= 2709)) || ((pixel_index >= 2713) && (pixel_index <= 2720)) || ((pixel_index >= 2724) && (pixel_index <= 2730)) || ((pixel_index >= 2733) && (pixel_index <= 2739)) || ((pixel_index >= 2742) && (pixel_index <= 2746)) || ((pixel_index >= 2749) && (pixel_index <= 2805)) || ((pixel_index >= 2809) && (pixel_index <= 2815)) || ((pixel_index >= 2819) && (pixel_index <= 2826)) || ((pixel_index >= 2830) && (pixel_index <= 2835)) || ((pixel_index >= 2838) && (pixel_index <= 2842)) || ((pixel_index >= 2845) && (pixel_index <= 2846)) || ((pixel_index >= 2856) && (pixel_index <= 2901)) || ((pixel_index >= 2914) && (pixel_index <= 2922)) || ((pixel_index >= 2928) && (pixel_index <= 2930)) || ((pixel_index >= 2933) && (pixel_index <= 2938)) || ((pixel_index >= 2954) && (pixel_index <= 2997)) || ((pixel_index >= 3012) && (pixel_index <= 3018)) || ((pixel_index >= 3021) && (pixel_index <= 3022)) || ((pixel_index >= 3028) && (pixel_index <= 3033)) || ((pixel_index >= 3039) && (pixel_index <= 3046)) || ((pixel_index >= 3051) && (pixel_index <= 3093)) || ((pixel_index >= 3097) && (pixel_index <= 3104)) || ((pixel_index >= 3109) && (pixel_index <= 3129)) || ((pixel_index >= 3133) && (pixel_index <= 3143)) || ((pixel_index >= 3147) && (pixel_index <= 3189)) || ((pixel_index >= 3193) && (pixel_index <= 3202)) || ((pixel_index >= 3206) && (pixel_index <= 3225)) || ((pixel_index >= 3229) && (pixel_index <= 3240)) || ((pixel_index >= 3243) && (pixel_index <= 3285)) || ((pixel_index >= 3289) && (pixel_index <= 3299)) || ((pixel_index >= 3303) && (pixel_index <= 3322)) || ((pixel_index >= 3325) && (pixel_index <= 3336)) || ((pixel_index >= 3340) && (pixel_index <= 3381)) || ((pixel_index >= 3385) && (pixel_index <= 3395)) || ((pixel_index >= 3399) && (pixel_index <= 3418)) || ((pixel_index >= 3421) && (pixel_index <= 3432)) || ((pixel_index >= 3436) && (pixel_index <= 3477)) || ((pixel_index >= 3481) && (pixel_index <= 3491)) || ((pixel_index >= 3495) && (pixel_index <= 3514)) || ((pixel_index >= 3517) && (pixel_index <= 3528)) || ((pixel_index >= 3532) && (pixel_index <= 3573)) || ((pixel_index >= 3577) && (pixel_index <= 3587)) || ((pixel_index >= 3591) && (pixel_index <= 3610)) || ((pixel_index >= 3614) && (pixel_index <= 3624)) || ((pixel_index >= 3628) && (pixel_index <= 3669)) || ((pixel_index >= 3673) && (pixel_index <= 3683)) || ((pixel_index >= 3687) && (pixel_index <= 3706)) || ((pixel_index >= 3710) && (pixel_index <= 3720)) || ((pixel_index >= 3724) && (pixel_index <= 3765)) || ((pixel_index >= 3769) && (pixel_index <= 3779)) || ((pixel_index >= 3783) && (pixel_index <= 3802)) || ((pixel_index >= 3806) && (pixel_index <= 3815)) || ((pixel_index >= 3819) && (pixel_index <= 3861)) || ((pixel_index >= 3865) && (pixel_index <= 3874)) || ((pixel_index >= 3878) && (pixel_index <= 3899)) || ((pixel_index >= 3903) && (pixel_index <= 3911)) || ((pixel_index >= 3915) && (pixel_index <= 3957)) || ((pixel_index >= 3961) && (pixel_index <= 3969)) || ((pixel_index >= 3974) && (pixel_index <= 3995)) || ((pixel_index >= 3999) && (pixel_index <= 4006)) || ((pixel_index >= 4010) && (pixel_index <= 4053)) || ((pixel_index >= 4057) && (pixel_index <= 4063)) || ((pixel_index >= 4069) && (pixel_index <= 4092)) || ((pixel_index >= 4097) && (pixel_index <= 4101)) || ((pixel_index >= 4106) && (pixel_index <= 4149)) || ((pixel_index >= 4164) && (pixel_index <= 4189)) || ((pixel_index >= 4201) && (pixel_index <= 4246)) || ((pixel_index >= 4258) && (pixel_index <= 4286)) || (pixel_index >= 4295) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 1291 || pixel_index == 1387 || pixel_index == 1483 || pixel_index == 1579 || pixel_index == 1675 || pixel_index == 1771 || pixel_index == 1867 || pixel_index == 1963 || pixel_index == 1965 || pixel_index == 2059 || pixel_index == 2155 || pixel_index == 2251 || pixel_index == 2347 || pixel_index == 2358 || pixel_index == 2443 || pixel_index == 2539 || pixel_index == 2635 || pixel_index == 2731 || pixel_index == 2827 || pixel_index == 2923 || pixel_index == 3019 || pixel_index == 3034 || pixel_index == 3226 || pixel_index == 3816 || pixel_index == 4200) oled_data = 16'b1010010100010100;
    else if (pixel_index == 2049 || pixel_index == 2242 || pixel_index == 3130) oled_data = 16'b0101001010001010;
    else oled_data = 0;
    end
    
    else if (freq>=1975 && freq<2093) //B6
    begin 
    if (((pixel_index >= 0) && (pixel_index <= 1757)) || ((pixel_index >= 1769) && (pixel_index <= 1784)) || ((pixel_index >= 1795) && (pixel_index <= 1853)) || ((pixel_index >= 1867) && (pixel_index <= 1879)) || ((pixel_index >= 1891) && (pixel_index <= 1949)) || ((pixel_index >= 1952) && (pixel_index <= 1958)) || ((pixel_index >= 1964) && (pixel_index <= 1974)) || ((pixel_index >= 1978) && (pixel_index <= 1985)) || ((pixel_index >= 1987) && (pixel_index <= 2045)) || ((pixel_index >= 2048) && (pixel_index <= 2056)) || ((pixel_index >= 2060) && (pixel_index <= 2069)) || ((pixel_index >= 2073) && (pixel_index <= 2141)) || ((pixel_index >= 2144) && (pixel_index <= 2153)) || ((pixel_index >= 2157) && (pixel_index <= 2164)) || ((pixel_index >= 2168) && (pixel_index <= 2237)) || ((pixel_index >= 2240) && (pixel_index <= 2249)) || ((pixel_index >= 2253) && (pixel_index <= 2260)) || ((pixel_index >= 2263) && (pixel_index <= 2333)) || ((pixel_index >= 2336) && (pixel_index <= 2345)) || ((pixel_index >= 2349) && (pixel_index <= 2355)) || ((pixel_index >= 2359) && (pixel_index <= 2429)) || ((pixel_index >= 2432) && (pixel_index <= 2441)) || ((pixel_index >= 2445) && (pixel_index <= 2451)) || ((pixel_index >= 2455) && (pixel_index <= 2525)) || ((pixel_index >= 2528) && (pixel_index <= 2537)) || ((pixel_index >= 2541) && (pixel_index <= 2547)) || ((pixel_index >= 2550) && (pixel_index <= 2621)) || ((pixel_index >= 2624) && (pixel_index <= 2632)) || ((pixel_index >= 2636) && (pixel_index <= 2642)) || ((pixel_index >= 2646) && (pixel_index <= 2717)) || ((pixel_index >= 2720) && (pixel_index <= 2728)) || ((pixel_index >= 2732) && (pixel_index <= 2738)) || ((pixel_index >= 2742) && (pixel_index <= 2813)) || ((pixel_index >= 2816) && (pixel_index <= 2822)) || ((pixel_index >= 2827) && (pixel_index <= 2834)) || pixel_index == 2838 || ((pixel_index >= 2849) && (pixel_index <= 2909)) || ((pixel_index >= 2921) && (pixel_index <= 2930)) || ((pixel_index >= 2946) && (pixel_index <= 3005)) || ((pixel_index >= 3020) && (pixel_index <= 3026)) || ((pixel_index >= 3032) && (pixel_index <= 3039)) || ((pixel_index >= 3043) && (pixel_index <= 3101)) || ((pixel_index >= 3104) && (pixel_index <= 3111)) || ((pixel_index >= 3117) && (pixel_index <= 3122)) || ((pixel_index >= 3126) && (pixel_index <= 3136)) || ((pixel_index >= 3140) && (pixel_index <= 3197)) || ((pixel_index >= 3200) && (pixel_index <= 3209)) || ((pixel_index >= 3214) && (pixel_index <= 3218)) || ((pixel_index >= 3222) && (pixel_index <= 3232)) || ((pixel_index >= 3236) && (pixel_index <= 3293)) || ((pixel_index >= 3296) && (pixel_index <= 3306)) || ((pixel_index >= 3310) && (pixel_index <= 3314)) || ((pixel_index >= 3318) && (pixel_index <= 3328)) || ((pixel_index >= 3332) && (pixel_index <= 3389)) || ((pixel_index >= 3392) && (pixel_index <= 3402)) || ((pixel_index >= 3406) && (pixel_index <= 3410)) || ((pixel_index >= 3414) && (pixel_index <= 3425)) || ((pixel_index >= 3428) && (pixel_index <= 3485)) || ((pixel_index >= 3488) && (pixel_index <= 3499)) || ((pixel_index >= 3503) && (pixel_index <= 3506)) || ((pixel_index >= 3510) && (pixel_index <= 3521)) || ((pixel_index >= 3524) && (pixel_index <= 3581)) || ((pixel_index >= 3584) && (pixel_index <= 3595)) || ((pixel_index >= 3599) && (pixel_index <= 3602)) || ((pixel_index >= 3606) && (pixel_index <= 3617)) || ((pixel_index >= 3620) && (pixel_index <= 3677)) || ((pixel_index >= 3680) && (pixel_index <= 3691)) || ((pixel_index >= 3694) && (pixel_index <= 3699)) || ((pixel_index >= 3702) && (pixel_index <= 3712)) || ((pixel_index >= 3716) && (pixel_index <= 3773)) || ((pixel_index >= 3776) && (pixel_index <= 3786)) || ((pixel_index >= 3790) && (pixel_index <= 3795)) || ((pixel_index >= 3799) && (pixel_index <= 3808)) || ((pixel_index >= 3812) && (pixel_index <= 3869)) || ((pixel_index >= 3872) && (pixel_index <= 3882)) || ((pixel_index >= 3886) && (pixel_index <= 3891)) || ((pixel_index >= 3895) && (pixel_index <= 3904)) || ((pixel_index >= 3908) && (pixel_index <= 3965)) || ((pixel_index >= 3968) && (pixel_index <= 3977)) || ((pixel_index >= 3981) && (pixel_index <= 3988)) || ((pixel_index >= 3992) && (pixel_index <= 3999)) || ((pixel_index >= 4003) && (pixel_index <= 4061)) || ((pixel_index >= 4064) && (pixel_index <= 4070)) || ((pixel_index >= 4077) && (pixel_index <= 4084)) || ((pixel_index >= 4089) && (pixel_index <= 4093)) || ((pixel_index >= 4098) && (pixel_index <= 4157)) || ((pixel_index >= 4171) && (pixel_index <= 4181)) || ((pixel_index >= 4193) && (pixel_index <= 4253)) || ((pixel_index >= 4265) && (pixel_index <= 4279)) || (pixel_index >= 4287) && (pixel_index <= 6143)) oled_data = 16'b1111011110011110;
    else if (pixel_index == 2156 || pixel_index == 3403 || pixel_index == 3598) oled_data = 16'b0101001010001010;
    else if (pixel_index == 2454) oled_data = 16'b0101010100001010;
    else if (pixel_index == 2839 || pixel_index == 3213 || pixel_index == 3329 || pixel_index == 3502 || pixel_index == 3907) oled_data = 16'b1010010100010100;
    else oled_data = 0;
    end
 
    
    
    end
    
    
endmodule


